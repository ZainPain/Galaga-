��S p r i t e T a b l e B   =   ' { ' { 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 } ,  
 ' { 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h d e , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 } ,  
 ' { 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h d e , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 } ,  
 ' { 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h d e , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 } ,  
 ' { 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 } ,  
 ' { 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 } ,  
 ' { 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 } ,  
 ' { 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 } ,  
 ' { 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h d e , 8 ' h 0 , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h 0 , 8 ' h d e , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 } ,  
 ' { 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h 0 , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 } ,  
 ' { 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 } ,  
 ' { 8 ' h 0 , 8 ' h d e , 8 ' h 0 , 8 ' h 0 , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h 0 , 8 ' h d e , 8 ' h 0 , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h 0 , 8 ' h 0 , 8 ' h d e , 8 ' h 0 } ,  
 ' { 8 ' h 0 , 8 ' h d e , 8 ' h 0 , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h 0 , 8 ' h d e , 8 ' h 0 } ,  
 ' { 8 ' h 0 , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h 0 , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h 0 , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h 0 } ,  
 ' { 8 ' h 0 , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h d e , 8 ' h d e , 8 ' h d e , 8 ' h 0 } ,  
 ' { 8 ' h 0 , 8 ' h d e , 8 ' h d e , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h d e , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h d e , 8 ' h d e , 8 ' h 0 } ,  
 ' { 8 ' h 0 , 8 ' h d e , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h d e , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h d e , 8 ' h 0 } ,  
 ' { 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 } ,  
 ' { 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 , 8 ' h 0 } } ;  
 