/* This is a Constant Array in Hardware which is utilized for the GalagaLogo */
module GalagaLogo(input [9:0] SpriteX, SpriteY,
            output [7:0] SpriteR, SpriteG, SpriteB);

parameter bit [7:0] SpriteTableR[111:0][226:0] = '{'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h25,8'h24,8'h24,8'h23,8'h23,8'h22,8'h22,8'h22,8'h22,8'h22,8'h22,8'h22,8'h22,8'h22,8'h22,8'h22,8'h22,8'h22,8'h23,8'h23,8'h23,8'h24,8'h24,8'h24,8'h25,8'h25,8'h25,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h25,8'h25,8'h25,8'h2b,8'h32,8'h3b,8'h43,8'h52,8'h5b,8'h63,8'h6f,8'h77,8'h7a,8'h7c,8'h7b,8'h7a,8'h7c,8'h7b,8'h7c,8'h7e,8'h7e,8'h7e,8'h7a,8'h73,8'h70,8'h6d,8'h66,8'h60,8'h5b,8'h54,8'h4c,8'h45,8'h37,8'h32,8'h2e,8'h27,8'h25,8'h25,8'h25,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h28,8'h2b,8'h33,8'h48,8'h4d,8'h4e,8'h50,8'h6b,8'h92,8'haa,8'hbc,8'hc5,8'hda,8'he5,8'hed,8'hf6,8'hfc,8'hff,8'hff,8'hfd,8'hfb,8'hfe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hfb,8'hf5,8'hf3,8'hf4,8'hee,8'hea,8'he5,8'he1,8'hd5,8'hc9,8'hba,8'hb5,8'h94,8'h5c,8'h4b,8'h4b,8'h4b,8'h48,8'h40,8'h2d,8'h29,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h25,8'h00,8'h2b,8'h33,8'h3d,8'h4e,8'h6a,8'h8c,8'haa,8'hc1,8'hde,8'he6,8'he8,8'heb,8'hf5,8'hfd,8'hff,8'hff,8'hff,8'hf8,8'hf1,8'he9,8'he0,8'hd2,8'hcb,8'hc4,8'hbe,8'hb4,8'ha9,8'ha9,8'ha3,8'ha1,8'ha1,8'ha1,8'ha4,8'hb4,8'hbb,8'hbf,8'hc6,8'hcf,8'hd5,8'he0,8'hee,8'hf5,8'hfa,8'hff,8'hfc,8'hf0,8'hea,8'he6,8'he6,8'hdf,8'hcd,8'hb0,8'h98,8'h75,8'h51,8'h41,8'h35,8'h2c,8'h28,8'h25,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h24,8'h25,8'h2b,8'h38,8'h4a,8'h69,8'h8e,8'hb4,8'hd0,8'he4,8'hf2,8'hfd,8'hff,8'hff,8'hff,8'hfd,8'hf1,8'he2,8'hcf,8'hba,8'ha5,8'h96,8'h80,8'h6d,8'h60,8'h50,8'h4d,8'h44,8'h39,8'h3b,8'h42,8'h42,8'h3c,8'h3f,8'h3e,8'h41,8'h43,8'h42,8'h40,8'h43,8'h42,8'h38,8'h36,8'h38,8'h43,8'h47,8'h58,8'h63,8'h67,8'h79,8'h96,8'had,8'hc7,8'hdd,8'hed,8'hfc,8'hff,8'hff,8'hff,8'hfa,8'he8,8'hd8,8'hb8,8'h94,8'h75,8'h52,8'h3f,8'h2e,8'h26,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h2f,8'h50,8'h6c,8'h8d,8'hb5,8'hd6,8'hf1,8'hff,8'hff,8'hff,8'hff,8'hf2,8'he1,8'hcc,8'haf,8'h8d,8'h76,8'h62,8'h4f,8'h45,8'h44,8'h42,8'h46,8'h47,8'h4e,8'h53,8'h5b,8'h5f,8'h62,8'h61,8'h65,8'h65,8'h66,8'h62,8'h63,8'h69,8'h69,8'h69,8'h64,8'h63,8'h60,8'h64,8'h5e,8'h5e,8'h5c,8'h61,8'h5c,8'h50,8'h4a,8'h49,8'h48,8'h42,8'h41,8'h43,8'h4e,8'h62,8'h72,8'h8d,8'hae,8'hc6,8'hdc,8'hef,8'hff,8'hff,8'hff,8'hf7,8'he1,8'hc0,8'h93,8'h6c,8'h44,8'h28,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h00,8'h27,8'h30,8'h49,8'h6c,8'h9d,8'hd3,8'hed,8'hfd,8'hff,8'hff,8'hff,8'hea,8'hcd,8'ha4,8'h81,8'h5c,8'h4d,8'h46,8'h46,8'h4a,8'h51,8'h55,8'h57,8'h60,8'h68,8'h70,8'h70,8'h71,8'h6c,8'h69,8'h6d,8'h62,8'h64,8'h66,8'h61,8'h60,8'h62,8'h5f,8'h59,8'h5f,8'h5d,8'h5a,8'h52,8'h55,8'h58,8'h5b,8'h5e,8'h5c,8'h5f,8'h68,8'h63,8'h6a,8'h72,8'h6f,8'h71,8'h6b,8'h69,8'h5e,8'h53,8'h50,8'h4d,8'h4e,8'h49,8'h49,8'h50,8'h5e,8'h77,8'ha3,8'hc9,8'he7,8'hfe,8'hff,8'hfd,8'hec,8'hc9,8'h94,8'h71,8'h4a,8'h2f,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h28,8'h2a,8'h32,8'h48,8'h76,8'haf,8'hd8,8'hef,8'hfd,8'hff,8'hff,8'hf5,8'hdc,8'hb3,8'h80,8'h50,8'h43,8'h44,8'h4f,8'h5c,8'h66,8'h67,8'h6d,8'h7b,8'h7b,8'h7a,8'h76,8'h6d,8'h69,8'h63,8'h5c,8'h63,8'h5b,8'h4f,8'h49,8'h41,8'h3d,8'h3b,8'h41,8'h41,8'h40,8'h43,8'h43,8'h40,8'h41,8'h42,8'h40,8'h40,8'h3e,8'h3e,8'h40,8'h44,8'h43,8'h42,8'h35,8'h3f,8'h46,8'h3e,8'h43,8'h55,8'h60,8'h5e,8'h62,8'h65,8'h6c,8'h74,8'h65,8'h61,8'h5a,8'h52,8'h4a,8'h4d,8'h44,8'h4f,8'h76,8'ha2,8'hcb,8'hed,8'hfd,8'hf9,8'hea,8'hdb,8'hac,8'h68,8'h46,8'h30,8'h26,8'h25,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h29,8'h36,8'h54,8'h7a,8'h8f,8'hb9,8'he0,8'hfa,8'hfc,8'hf0,8'hda,8'had,8'h96,8'h93,8'h7d,8'h6b,8'h54,8'h4b,8'h5c,8'h75,8'h81,8'h8a,8'h85,8'h72,8'h64,8'h5d,8'h5b,8'h4d,8'h4f,8'h5a,8'h63,8'h69,8'h6c,8'h79,8'h8a,8'h91,8'h8f,8'h8d,8'h8d,8'h8b,8'h8e,8'ha5,8'hb2,8'hbe,8'hc8,8'hcf,8'hd0,8'hcf,8'hd0,8'hd2,8'hd3,8'hd2,8'hd2,8'hd3,8'hd0,8'hc4,8'hb7,8'ha3,8'h97,8'h8b,8'h84,8'h8b,8'h91,8'h96,8'h8d,8'h76,8'h63,8'h63,8'h5d,8'h54,8'h4e,8'h4f,8'h56,8'h62,8'h65,8'h5e,8'h60,8'h4b,8'h4d,8'h58,8'h6a,8'h82,8'h92,8'ha5,8'hd1,8'hec,8'hef,8'he1,8'h91,8'h2d,8'h31,8'h46,8'h30,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h27,8'h3b,8'h74,8'hae,8'hdc,8'hf8,8'hff,8'hff,8'hf7,8'hd8,8'h9e,8'h70,8'h54,8'h45,8'h4b,8'h61,8'h6e,8'h78,8'h7e,8'h80,8'h7d,8'h75,8'h6a,8'h62,8'h4f,8'h40,8'h43,8'h49,8'h57,8'h6c,8'h87,8'ha8,8'hc8,8'he2,8'hef,8'hf8,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfe,8'hfd,8'hfb,8'hff,8'hff,8'hfd,8'hfe,8'hfc,8'hfd,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hf7,8'hec,8'hde,8'hc5,8'haa,8'h8d,8'h73,8'h5e,8'h4f,8'h47,8'h44,8'h4f,8'h5f,8'h6a,8'h6b,8'h65,8'h55,8'h49,8'h41,8'h45,8'h65,8'h9b,8'hcc,8'h8b,8'h44,8'ha3,8'hd5,8'h9c,8'h5c,8'h30,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h2e,8'h4b,8'h80,8'hb4,8'he5,8'hfd,8'hfa,8'hf3,8'hd9,8'had,8'h75,8'h52,8'h4b,8'h59,8'h6b,8'h7d,8'h80,8'h7b,8'h74,8'h74,8'h67,8'h5f,8'h58,8'h48,8'h44,8'h56,8'h6c,8'h8c,8'hb3,8'hd6,8'hea,8'hfb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfa,8'hf2,8'hee,8'hed,8'he8,8'he7,8'he5,8'hdf,8'hcf,8'hc8,8'hc2,8'hcd,8'hb5,8'hb2,8'ha9,8'hab,8'ha8,8'ha1,8'hb1,8'hc2,8'hb7,8'hb0,8'hbb,8'hca,8'hd5,8'hdf,8'he5,8'he8,8'hec,8'hed,8'hef,8'hf0,8'hf4,8'hfb,8'hff,8'hff,8'hff,8'hff,8'hf8,8'hea,8'hd7,8'hb7,8'h8f,8'h72,8'h56,8'h49,8'h4c,8'h5d,8'h63,8'h6a,8'h6d,8'h60,8'h4b,8'h38,8'h36,8'h27,8'h5d,8'hd8,8'hf8,8'hf6,8'he0,8'ha4,8'h66,8'h3f,8'h2a,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h28,8'h29,8'h31,8'h40,8'h43,8'h50,8'h66,8'h67,8'h54,8'h43,8'h33,8'h29,8'h27,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h2c,8'h41,8'h6e,8'hab,8'hdb,8'hf4,8'hfb,8'he8,8'hbc,8'h7d,8'h68,8'h64,8'h5e,8'h5d,8'h64,8'h70,8'h7c,8'h7a,8'h6e,8'h5b,8'h4a,8'h44,8'h5a,8'h72,8'h94,8'hb8,8'hc5,8'hca,8'he6,8'hf5,8'hff,8'hff,8'hff,8'hff,8'hfa,8'hef,8'he2,8'hcc,8'hb0,8'h96,8'h83,8'h72,8'h62,8'h5c,8'h58,8'h53,8'h50,8'h4b,8'h43,8'h3d,8'h3c,8'h47,8'h31,8'h37,8'h33,8'h28,8'h3a,8'h34,8'h31,8'h43,8'h3b,8'h2b,8'h3c,8'h42,8'h4a,8'h49,8'h60,8'h5c,8'h58,8'h5e,8'h5a,8'h57,8'h60,8'h75,8'h8e,8'hab,8'hce,8'hdf,8'heb,8'hf7,8'hff,8'hff,8'hfa,8'hf5,8'he3,8'hca,8'hc2,8'hb7,8'h91,8'h6d,8'h56,8'h47,8'h4e,8'h44,8'h27,8'h40,8'h71,8'h7c,8'h70,8'h86,8'hc9,8'hea,8'hee,8'hd7,8'ha9,8'h7a,8'h43,8'h2b,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h00,8'h2c,8'h3a,8'h54,8'h77,8'h9f,8'hab,8'hc2,8'hd9,8'he3,8'heb,8'hf4,8'hf5,8'hec,8'hdf,8'hc3,8'h9a,8'h56,8'h28,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h30,8'h4f,8'h91,8'hce,8'hef,8'hff,8'hfd,8'hdd,8'h92,8'h53,8'h3f,8'h45,8'h63,8'h6e,8'h66,8'h6e,8'h6a,8'h65,8'h5d,8'h49,8'h3a,8'h49,8'h70,8'ha3,8'hd7,8'hf2,8'hff,8'hff,8'hff,8'hff,8'hff,8'hf9,8'hec,8'hdf,8'hc8,8'ha8,8'h8b,8'h6c,8'h4e,8'h39,8'h2b,8'h23,8'h18,8'h11,8'h19,8'h1b,8'h15,8'h18,8'h12,8'h11,8'h24,8'h21,8'h1a,8'h12,8'h0a,8'h3d,8'h39,8'h21,8'h4a,8'h3b,8'h29,8'h27,8'h3d,8'h29,8'h1a,8'h19,8'h16,8'h23,8'h42,8'h38,8'h24,8'h1d,8'h17,8'h17,8'h1e,8'h15,8'h1c,8'h21,8'h2c,8'h45,8'h5f,8'h6f,8'h94,8'hbf,8'hd6,8'heb,8'hf6,8'hfb,8'hff,8'hff,8'hff,8'hf3,8'hd1,8'h6d,8'h31,8'h49,8'h32,8'h49,8'h61,8'h68,8'h5e,8'h52,8'h52,8'h6a,8'haa,8'he4,8'hfc,8'hf6,8'hcf,8'h88,8'h4a,8'h2d,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h2a,8'h3f,8'h61,8'h95,8'hc9,8'hec,8'hfb,8'hfe,8'hf6,8'heb,8'he0,8'hd0,8'hc8,8'hc9,8'hca,8'hcf,8'he4,8'hfe,8'hfa,8'hc0,8'h45,8'h25},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h27,8'h35,8'h50,8'h97,8'hd7,8'hf7,8'hf1,8'hdc,8'hc8,8'h91,8'h5c,8'h47,8'h52,8'h69,8'h76,8'h77,8'h6d,8'h5b,8'h54,8'h5f,8'h5e,8'h58,8'h78,8'haa,8'hd6,8'hf7,8'hff,8'hff,8'hfe,8'hf5,8'he3,8'hd5,8'hcf,8'hc1,8'had,8'h8a,8'h59,8'h43,8'h46,8'h4f,8'h5b,8'h60,8'h4c,8'h2e,8'h1b,8'h1f,8'h17,8'h16,8'h13,8'h0b,8'h12,8'h0c,8'h0a,8'h20,8'h2a,8'h2d,8'h27,8'h23,8'h1d,8'h0e,8'h18,8'h22,8'h19,8'h2e,8'h23,8'h30,8'h24,8'h21,8'h28,8'h3b,8'h6f,8'hb3,8'h98,8'h48,8'h27,8'h21,8'h20,8'h24,8'h28,8'h23,8'h13,8'h10,8'h2c,8'h25,8'h17,8'h18,8'h2a,8'h42,8'h6a,8'h99,8'hbc,8'hca,8'hd3,8'hdc,8'hed,8'hd5,8'h83,8'h66,8'h75,8'h8b,8'h6d,8'h58,8'h6c,8'h67,8'h66,8'h61,8'h57,8'h52,8'h69,8'ha9,8'hd5,8'he4,8'hee,8'hd2,8'h80,8'h3e,8'h33,8'h27,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h2e,8'h3f,8'h79,8'hc5,8'he7,8'hec,8'hdf,8'hd6,8'hc1,8'h9d,8'h80,8'h6a,8'h57,8'h45,8'h3c,8'h3b,8'h40,8'h44,8'h59,8'hb0,8'hfe,8'hf2,8'h88,8'h2c},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h29,8'h41,8'h76,8'hb5,8'hd9,8'hfa,8'hfc,8'hce,8'h7d,8'h58,8'h64,8'h5e,8'h68,8'h6f,8'h79,8'h70,8'h5b,8'h47,8'h3e,8'h4d,8'h82,8'hbc,8'hda,8'he6,8'hf6,8'hff,8'hff,8'hf8,8'hed,8'hcf,8'ha4,8'h7a,8'h54,8'h54,8'h6e,8'h40,8'h30,8'h32,8'h41,8'h7c,8'hb9,8'hd8,8'he4,8'he6,8'hd6,8'h92,8'h2f,8'h0f,8'h18,8'h18,8'h11,8'h12,8'h11,8'h0f,8'h0f,8'h13,8'h21,8'h25,8'h25,8'h24,8'h03,8'h0e,8'h1d,8'h26,8'h0e,8'h20,8'h23,8'h36,8'h15,8'h17,8'h28,8'h3b,8'h85,8'he9,8'hb6,8'h45,8'h24,8'h08,8'h10,8'h23,8'h2d,8'h34,8'h1e,8'h1d,8'h26,8'h18,8'h18,8'h07,8'h20,8'h1f,8'h29,8'h37,8'h50,8'h42,8'h47,8'h4a,8'h61,8'h7e,8'h85,8'h65,8'hbe,8'hfc,8'hf3,8'he2,8'hdc,8'hbf,8'h8a,8'h51,8'h49,8'h58,8'h62,8'h71,8'h70,8'h66,8'h8a,8'hcb,8'he6,8'hd0,8'hb7,8'h72,8'h3b,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h29,8'h3f,8'h67,8'ha8,8'hd0,8'hec,8'hde,8'h9e,8'h66,8'h4c,8'h4f,8'h58,8'h5b,8'h62,8'h64,8'h6d,8'h70,8'h71,8'h76,8'h76,8'h70,8'h58,8'h4e,8'hd5,8'hff,8'hc5,8'h34},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h27,8'h36,8'h70,8'hc6,8'hed,8'hfc,8'hf8,8'hc7,8'h76,8'h4c,8'h4e,8'h64,8'h77,8'h7d,8'h7f,8'h73,8'h66,8'h41,8'h39,8'h61,8'ha2,8'hd8,8'hf8,8'hff,8'hff,8'hff,8'hf8,8'he7,8'hd2,8'hb2,8'h80,8'h51,8'h2c,8'h24,8'h18,8'h24,8'h26,8'h1d,8'h47,8'h88,8'hc8,8'hec,8'hf9,8'hfd,8'hfe,8'hff,8'hf9,8'hd9,8'h5e,8'h17,8'h16,8'h13,8'h0c,8'h0d,8'h10,8'h0b,8'h10,8'h18,8'h21,8'h14,8'h16,8'h13,8'h0b,8'h15,8'h19,8'h20,8'h12,8'h1e,8'h20,8'h29,8'h13,8'h17,8'h10,8'h0c,8'h3f,8'h8b,8'h66,8'h2d,8'h0a,8'h14,8'h19,8'h08,8'h17,8'h25,8'h14,8'h1f,8'h15,8'h1c,8'h36,8'h19,8'h3f,8'h3d,8'h1a,8'h1d,8'h23,8'h1d,8'h3e,8'h2a,8'h41,8'h9f,8'h64,8'h41,8'h77,8'hb8,8'he2,8'hfa,8'hff,8'hff,8'hf7,8'hd6,8'h9e,8'h6a,8'h48,8'h4e,8'h61,8'h65,8'h57,8'h54,8'h83,8'hd2,8'hfd,8'hf0,8'hbb,8'h67,8'h37,8'h29,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h29,8'h3b,8'h73,8'hc6,8'hf0,8'hf0,8'hc3,8'h7b,8'h47,8'h39,8'h4f,8'h66,8'h6b,8'h66,8'h56,8'h4d,8'h4a,8'h65,8'h85,8'h83,8'h84,8'h86,8'h8d,8'h73,8'h3a,8'hc4,8'hff,8'hca,8'h35},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h25,8'h25,8'h25,8'h24,8'h25,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h39,8'h6d,8'hb1,8'hee,8'hf9,8'hdc,8'hb4,8'h89,8'h51,8'h50,8'h77,8'h82,8'h80,8'h6f,8'h60,8'h5c,8'h58,8'h62,8'h76,8'hbc,8'hf0,8'hff,8'hff,8'hf9,8'he3,8'hcb,8'hb2,8'h9e,8'h75,8'h57,8'h48,8'h2b,8'h23,8'h13,8'h19,8'h1c,8'h35,8'h58,8'h89,8'hd1,8'hf6,8'hfd,8'hf2,8'hd3,8'hb3,8'hb9,8'he2,8'hff,8'hf4,8'h89,8'h22,8'h1d,8'h1f,8'h20,8'h12,8'h10,8'h0c,8'h04,8'h0e,8'h18,8'h1c,8'h1d,8'h19,8'h15,8'h1c,8'h1f,8'h17,8'h16,8'h0f,8'h12,8'h12,8'h17,8'h16,8'h09,8'h08,8'h10,8'h3e,8'h27,8'h25,8'h1c,8'h21,8'h18,8'h12,8'h26,8'h22,8'h0f,8'h12,8'h11,8'h23,8'h3b,8'h1d,8'h31,8'h34,8'h10,8'h21,8'h27,8'h1f,8'h23,8'h4c,8'h9a,8'h72,8'h26,8'h25,8'h16,8'h28,8'h47,8'h77,8'ha8,8'hc2,8'hdd,8'hfa,8'hff,8'hee,8'hb7,8'h7b,8'h70,8'h6b,8'h62,8'h54,8'h4f,8'h64,8'h8f,8'hbc,8'he1,8'hea,8'hc2,8'h84,8'h50,8'h2b,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h2d,8'h58,8'h84,8'hc4,8'he3,8'hcd,8'haf,8'h7c,8'h47,8'h41,8'h5b,8'h65,8'h66,8'h6e,8'h72,8'h76,8'h6f,8'h66,8'h57,8'h38,8'h71,8'h86,8'h88,8'h8b,8'h85,8'h58,8'h5a,8'he8,8'hfa,8'h9e,8'h2f},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h25,8'h28,8'h31,8'h42,8'h45,8'h47,8'h52,8'h5a,8'h47,8'h3f,8'h2c,8'h00,8'h25,8'h00,8'h00,8'h00,8'h00,8'h25,8'h31,8'h62,8'haf,8'hf1,8'hfe,8'he0,8'h91,8'h53,8'h4d,8'h6b,8'h7c,8'h83,8'h7e,8'h74,8'h57,8'h40,8'h4a,8'h7d,8'hc6,8'hf3,8'hff,8'hff,8'hfb,8'he8,8'hcd,8'h98,8'h62,8'h3d,8'h2a,8'h27,8'h21,8'h23,8'h24,8'h24,8'h1c,8'h22,8'h33,8'h6d,8'hb9,8'he7,8'hf7,8'hfe,8'hf7,8'hc9,8'h7f,8'h49,8'h3b,8'h3c,8'h74,8'hf9,8'hfe,8'ha1,8'h26,8'h29,8'h30,8'h40,8'h24,8'h15,8'h1f,8'h15,8'h15,8'h16,8'h16,8'h1a,8'h1d,8'h19,8'h1b,8'h1c,8'h12,8'h12,8'h0e,8'h10,8'h12,8'h11,8'h10,8'h14,8'h1a,8'h15,8'h29,8'h23,8'h12,8'h23,8'h26,8'h13,8'h1f,8'h26,8'h1c,8'h0d,8'h14,8'h14,8'h16,8'h25,8'h28,8'h23,8'h3b,8'h25,8'h38,8'h41,8'h1d,8'h50,8'hc5,8'h8c,8'h23,8'h10,8'h14,8'h19,8'h1a,8'h0e,8'h0f,8'h24,8'h2d,8'h4f,8'h86,8'hbd,8'he2,8'hf9,8'hfb,8'hf3,8'hce,8'h91,8'h5c,8'h4b,8'h5f,8'h61,8'h5a,8'h66,8'ha0,8'he6,8'hfe,8'hdb,8'h81,8'h3d,8'h00,8'h00,8'h00,8'h25,8'h27,8'h43,8'h88,8'he3,8'hf2,8'hc1,8'h71,8'h46,8'h54,8'h6e,8'h78,8'h6e,8'h51,8'h54,8'h7d,8'hbb,8'he4,8'hf8,8'hf8,8'hf6,8'hdf,8'h52,8'h68,8'h89,8'h84,8'h87,8'h6e,8'h3c,8'ha5,8'hff,8'hcd,8'h4a,8'h25},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h28,8'h2b,8'h3d,8'h57,8'h72,8'h91,8'hae,8'hc8,8'hce,8'hd3,8'hdd,8'he1,8'hcf,8'hc1,8'h9c,8'h75,8'h59,8'h3b,8'h29,8'h28,8'h2e,8'h51,8'ha1,8'he1,8'hfe,8'hec,8'ha2,8'h59,8'h4b,8'h62,8'h76,8'h82,8'h76,8'h73,8'h63,8'h46,8'h4c,8'h84,8'hcd,8'hf9,8'hff,8'hfc,8'hf5,8'he3,8'hb7,8'h77,8'h43,8'h24,8'h12,8'h1b,8'h20,8'h21,8'h1c,8'h1a,8'h1f,8'h1a,8'h25,8'h60,8'haa,8'he5,8'hf9,8'hfb,8'hf4,8'hc4,8'h76,8'h43,8'h32,8'h49,8'h66,8'h49,8'h44,8'he6,8'hff,8'ha1,8'h25,8'h40,8'h41,8'h2d,8'h36,8'h3d,8'h21,8'h1f,8'h1a,8'h16,8'h16,8'h17,8'h15,8'h15,8'h18,8'h1d,8'h1a,8'h16,8'h12,8'h11,8'h11,8'h12,8'h11,8'h0d,8'h15,8'h13,8'h15,8'h14,8'h12,8'h1b,8'h1b,8'h17,8'h1d,8'h16,8'h08,8'h10,8'h19,8'h12,8'h12,8'h21,8'h1f,8'h1d,8'h22,8'h10,8'h20,8'h1d,8'h45,8'hc3,8'hba,8'h3a,8'h14,8'h1a,8'h1f,8'h18,8'h1c,8'h18,8'h13,8'h0c,8'h21,8'h4e,8'h36,8'h30,8'h5d,8'h99,8'hd6,8'hf2,8'hfe,8'hfc,8'he1,8'ha2,8'h6a,8'h55,8'h61,8'h5b,8'h4e,8'h66,8'haf,8'hf1,8'hef,8'hb1,8'h60,8'h2e,8'h28,8'h39,8'h7d,8'hc5,8'hef,8'hcf,8'h76,8'h47,8'h4c,8'h6f,8'h81,8'h7f,8'h65,8'h4f,8'h7a,8'hcd,8'hf6,8'hff,8'hfb,8'hf6,8'hf0,8'hf6,8'hde,8'h57,8'h6d,8'h89,8'h83,8'h87,8'h4e,8'h58,8'he8,8'hfd,8'h90,8'h2b,8'h25},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h00,8'h31,8'h57,8'h8c,8'haa,8'hc6,8'he0,8'hf0,8'hfb,8'hff,8'hff,8'hff,8'hff,8'hfa,8'hf8,8'hfd,8'hff,8'hff,8'hf8,8'he6,8'hc1,8'ha1,8'h9d,8'hb1,8'he1,8'hfa,8'hd4,8'h88,8'h6a,8'h5b,8'h67,8'h7c,8'h85,8'h7e,8'h68,8'h47,8'h51,8'h83,8'haa,8'hd5,8'hfa,8'hff,8'hf9,8'he1,8'hae,8'h77,8'h58,8'h30,8'h1d,8'h0e,8'h1b,8'h1d,8'h22,8'h21,8'h14,8'h12,8'h1f,8'h36,8'h71,8'ha8,8'he0,8'hf9,8'hfe,8'hdf,8'h98,8'h6d,8'h53,8'h4c,8'h5e,8'h64,8'h6b,8'h6b,8'h4c,8'h3c,8'he1,8'hff,8'ha8,8'h28,8'h2a,8'h29,8'h1d,8'h45,8'h60,8'h13,8'h13,8'h1b,8'h1e,8'h19,8'h1b,8'h18,8'h15,8'h15,8'h18,8'h18,8'h12,8'h11,8'h14,8'h12,8'h1f,8'h26,8'h28,8'h2c,8'h0b,8'h0b,8'h18,8'h24,8'h28,8'h11,8'h1f,8'h14,8'h13,8'h11,8'h15,8'h19,8'h12,8'h16,8'h0d,8'h18,8'h1b,8'h0f,8'h0b,8'h1f,8'h4f,8'hc3,8'hb9,8'h40,8'h20,8'h18,8'h2c,8'h3b,8'h1d,8'h1f,8'h19,8'h18,8'h20,8'h1f,8'h3b,8'h28,8'h1f,8'h24,8'h34,8'h5c,8'h71,8'h8c,8'hbd,8'hf4,8'hff,8'he6,8'hbe,8'h94,8'h68,8'h4f,8'h4d,8'h63,8'h6f,8'h96,8'hdd,8'hdf,8'haa,8'h9f,8'hc1,8'hdf,8'ha2,8'h6d,8'h5b,8'h54,8'h5f,8'h7e,8'h87,8'h61,8'h57,8'h8e,8'hc5,8'hf0,8'hfd,8'he8,8'hb1,8'h87,8'h7c,8'ha0,8'hef,8'ha4,8'h47,8'h78,8'h89,8'h89,8'h67,8'h4a,8'hbb,8'hff,8'hca,8'h4a,8'h25,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h2e,8'h56,8'ha8,8'he1,8'hf7,8'hff,8'hff,8'hff,8'hff,8'hf9,8'he6,8'hcd,8'had,8'h93,8'h7b,8'h74,8'h86,8'h9f,8'hc9,8'hea,8'hff,8'hff,8'hff,8'hff,8'hff,8'hf4,8'haf,8'h57,8'h46,8'h70,8'h85,8'h7b,8'h81,8'h74,8'h49,8'h3c,8'h65,8'hbd,8'hf9,8'hff,8'hff,8'hf4,8'he0,8'ha9,8'h5e,8'h2a,8'h14,8'h0e,8'h0d,8'h10,8'h1f,8'h20,8'h20,8'h24,8'h19,8'h0c,8'h25,8'h58,8'haf,8'hef,8'hff,8'hfe,8'heb,8'ha6,8'h4f,8'h3b,8'h56,8'h71,8'h6c,8'h68,8'h6c,8'h6e,8'h6e,8'h4e,8'h3e,8'he1,8'hfa,8'hcb,8'h40,8'h20,8'h1f,8'h1e,8'h24,8'h23,8'h17,8'h1f,8'h1b,8'h19,8'h15,8'h1b,8'h16,8'h12,8'h07,8'h0b,8'h13,8'h1a,8'h1e,8'h18,8'h16,8'h24,8'h33,8'h31,8'h27,8'h14,8'h0e,8'h12,8'h20,8'h22,8'h0f,8'h20,8'h14,8'h0e,8'h15,8'h16,8'h1a,8'h16,8'h19,8'h24,8'h14,8'h11,8'h14,8'h15,8'h50,8'hd1,8'hd4,8'h46,8'h14,8'h1c,8'h11,8'h44,8'h4e,8'h21,8'h1b,8'h1d,8'h1c,8'h1d,8'h1b,8'h14,8'h1d,8'h4b,8'h3f,8'h41,8'h46,8'h20,8'h23,8'h31,8'h6e,8'hb8,8'he8,8'hfd,8'hff,8'he4,8'h99,8'h5a,8'h50,8'h56,8'h4c,8'h63,8'ha8,8'hec,8'hf3,8'hc1,8'h63,8'h38,8'h51,8'h79,8'h78,8'h7c,8'h74,8'h52,8'h50,8'hb1,8'hfa,8'hfc,8'he3,8'ha5,8'h62,8'h36,8'h29,8'h2c,8'h8c,8'he6,8'h60,8'h59,8'h82,8'h84,8'h6d,8'h37,8'h81,8'hfa,8'hf2,8'h7e,8'h28,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h30,8'h57,8'h99,8'hd6,8'hf8,8'hff,8'hff,8'hf6,8'he7,8'hd6,8'haa,8'h80,8'h63,8'h55,8'h54,8'h5b,8'h5d,8'h5c,8'h5c,8'h4e,8'h50,8'h68,8'h96,8'hc3,8'he2,8'he4,8'hc0,8'h77,8'h4b,8'h63,8'h77,8'h80,8'h81,8'h6c,8'h64,8'h55,8'h62,8'hb1,8'hf2,8'hff,8'hfc,8'he8,8'hd8,8'hbe,8'h61,8'h29,8'h0d,8'h11,8'h16,8'h14,8'h21,8'h18,8'h25,8'h43,8'h29,8'h14,8'h26,8'h45,8'h83,8'hd8,8'hf8,8'hf6,8'he6,8'hb5,8'h5c,8'h34,8'h49,8'h62,8'h71,8'h72,8'h6c,8'h6a,8'h70,8'h6f,8'h6d,8'h4a,8'h3f,8'he1,8'hf7,8'haf,8'h2a,8'h1f,8'h22,8'h23,8'h1c,8'h0c,8'h1b,8'h1b,8'h18,8'h17,8'h21,8'h21,8'h1a,8'h28,8'h24,8'h15,8'h14,8'h1b,8'h11,8'h1a,8'h21,8'h22,8'h1f,8'h25,8'h29,8'h24,8'h14,8'h20,8'h22,8'h1d,8'h18,8'h1f,8'h16,8'h10,8'h10,8'h1a,8'h1e,8'h18,8'h0e,8'h13,8'h14,8'h1d,8'h25,8'h4b,8'hc4,8'he2,8'h6a,8'h17,8'h22,8'h2a,8'h4c,8'h90,8'h9b,8'h54,8'h24,8'h23,8'h2b,8'h22,8'h19,8'h1a,8'h11,8'h25,8'h25,8'h44,8'h2c,8'h36,8'h3b,8'h18,8'h1f,8'h4a,8'h75,8'hac,8'hdf,8'hf6,8'hfc,8'hd4,8'h86,8'h63,8'h65,8'h5b,8'h4c,8'h71,8'h7a,8'h47,8'h42,8'h65,8'h75,8'h73,8'h70,8'h6c,8'h5e,8'h6f,8'hc8,8'hfe,8'hec,8'hb9,8'h6b,8'h32,8'h27,8'h26,8'h26,8'h55,8'hd8,8'hbd,8'h44,8'h79,8'h85,8'h80,8'h4d,8'h5f,8'hdd,8'hfa,8'haf,8'h3c,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2e,8'h65,8'hae,8'hd9,8'hfb,8'hff,8'hff,8'hee,8'hb1,8'h6d,8'h62,8'h71,8'h6c,8'h68,8'h6c,8'h77,8'h82,8'h88,8'h86,8'h83,8'h84,8'h7e,8'h72,8'h6e,8'h65,8'h65,8'h6f,8'h58,8'h54,8'h5d,8'h6a,8'h7a,8'h77,8'h71,8'h57,8'h47,8'h7b,8'hc3,8'heb,8'hff,8'hfd,8'hee,8'hd3,8'h8f,8'h52,8'h42,8'h1f,8'h12,8'h21,8'h38,8'h23,8'h22,8'h22,8'h19,8'h23,8'h32,8'h24,8'h37,8'h8b,8'hd1,8'hf1,8'hfe,8'hff,8'hed,8'ha9,8'h74,8'h56,8'h62,8'h59,8'h4b,8'h76,8'h6d,8'h6a,8'h6b,8'h6d,8'h71,8'h6e,8'h48,8'h3f,8'he2,8'hf9,8'h98,8'h20,8'h1b,8'h11,8'h11,8'h14,8'h0f,8'h0f,8'h05,8'h19,8'h23,8'h32,8'h32,8'h1d,8'h20,8'h24,8'h1f,8'h1a,8'h1e,8'h22,8'h23,8'h23,8'h1d,8'h1f,8'h28,8'h1d,8'h15,8'h10,8'h13,8'h12,8'h15,8'h1d,8'h1b,8'h15,8'h13,8'h13,8'h1d,8'h20,8'h16,8'h04,8'h0f,8'h1d,8'h20,8'h5c,8'hce,8'he7,8'h75,8'h22,8'h10,8'h27,8'h52,8'h93,8'he4,8'hec,8'h96,8'h2e,8'h2b,8'h54,8'h2e,8'h11,8'h1d,8'h16,8'h0d,8'h1d,8'h27,8'h1f,8'h26,8'h2c,8'h1a,8'h22,8'h2e,8'h35,8'h3f,8'h49,8'h73,8'hbe,8'hf3,8'hf3,8'hd8,8'hb0,8'h6f,8'h49,8'h4e,8'h57,8'h64,8'h6d,8'h77,8'h75,8'h79,8'h60,8'h50,8'h9b,8'he7,8'hfa,8'hda,8'h78,8'h3f,8'h27,8'h25,8'h26,8'h25,8'h37,8'had,8'hdb,8'h61,8'h64,8'h87,8'h7f,8'h4c,8'h50,8'hcf,8'hf9,8'hbb,8'h46,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h27,8'h47,8'h90,8'hdf,8'hfa,8'hff,8'hff,8'hec,8'hb1,8'h66,8'h47,8'h5d,8'h74,8'h80,8'h81,8'h82,8'h7f,8'h6d,8'h61,8'h53,8'h47,8'h41,8'h3e,8'h6f,8'h8b,8'h83,8'h7e,8'h77,8'h71,8'h63,8'h71,8'h76,8'h75,8'h7e,8'h65,8'h40,8'h5b,8'hae,8'hf2,8'hff,8'hff,8'hf3,8'hd2,8'h83,8'h47,8'h2b,8'h11,8'h13,8'h19,8'h19,8'h24,8'h47,8'h21,8'h25,8'h22,8'h16,8'h19,8'h0a,8'h40,8'hc1,8'hf5,8'hff,8'hfe,8'hff,8'hff,8'hff,8'hf4,8'hf1,8'hf2,8'hf2,8'hc9,8'h4c,8'h5b,8'h75,8'h6e,8'h6f,8'h71,8'h71,8'h6e,8'h4b,8'h40,8'he2,8'hfa,8'h98,8'h22,8'h1a,8'h0e,8'h0e,8'h11,8'h13,8'h13,8'h0d,8'h0c,8'h1f,8'h2f,8'h52,8'h1f,8'h05,8'h1d,8'h28,8'h23,8'h26,8'h32,8'h25,8'h27,8'h16,8'h12,8'h0c,8'h00,8'h0c,8'h14,8'h0f,8'h10,8'h13,8'h17,8'h15,8'h14,8'h13,8'h0d,8'h0b,8'h0e,8'h07,8'h0e,8'h11,8'h17,8'h4c,8'hcc,8'hf7,8'h9c,8'h22,8'h18,8'h14,8'h1a,8'h24,8'h53,8'hd6,8'he0,8'h5f,8'h11,8'h1c,8'h26,8'h1a,8'h12,8'h21,8'h20,8'h18,8'h20,8'h25,8'h16,8'h0e,8'h12,8'h14,8'h19,8'h1d,8'h20,8'h0e,8'h06,8'h25,8'h3c,8'h84,8'hd7,8'hf5,8'hfd,8'he0,8'h94,8'h4e,8'h4d,8'h63,8'h6d,8'h7b,8'h7b,8'h72,8'h4c,8'ha1,8'hf7,8'hfc,8'he0,8'h6f,8'h2a,8'h25,8'h26,8'h26,8'h26,8'h28,8'h78,8'hef,8'h95,8'h42,8'h83,8'h8c,8'h65,8'h44,8'hb4,8'hff,8'hde,8'h5f,8'h25,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h2e,8'h60,8'hc1,8'hf5,8'hff,8'hff,8'hdf,8'hbd,8'h7c,8'h4e,8'h60,8'h7c,8'h84,8'h75,8'h69,8'h66,8'h6b,8'h72,8'h5c,8'h63,8'h85,8'h9c,8'h89,8'h48,8'h69,8'h86,8'h81,8'h81,8'h84,8'h7a,8'h74,8'h74,8'h78,8'h66,8'h5f,8'h62,8'h8e,8'he4,8'hff,8'hff,8'hec,8'hce,8'h94,8'h4f,8'h26,8'h1a,8'h1b,8'h12,8'h1a,8'h18,8'h19,8'h20,8'h0f,8'h10,8'h31,8'h30,8'h34,8'h27,8'h26,8'h57,8'hd8,8'hee,8'hf0,8'hf0,8'hee,8'hee,8'hf0,8'hf5,8'hf6,8'hf8,8'hfb,8'hf9,8'h75,8'h4b,8'h73,8'h71,8'h71,8'h6e,8'h6a,8'h6b,8'h4e,8'h40,8'he3,8'hfb,8'h96,8'h21,8'h1d,8'h17,8'h11,8'h13,8'h17,8'h19,8'h1d,8'h26,8'h31,8'h2f,8'h29,8'h18,8'h1f,8'h15,8'h04,8'h1f,8'h29,8'h1c,8'h21,8'h1e,8'h0b,8'h0d,8'h10,8'h0b,8'h09,8'h13,8'h10,8'h18,8'h19,8'h18,8'h19,8'h11,8'h0a,8'h05,8'h0a,8'h0b,8'h05,8'h1f,8'h24,8'h53,8'hc9,8'hf4,8'hbd,8'h3a,8'h16,8'h1d,8'h16,8'h1d,8'h20,8'h2f,8'h74,8'h7f,8'h2a,8'h20,8'h18,8'h1f,8'h20,8'h20,8'h13,8'h1f,8'h30,8'h20,8'h2e,8'h23,8'h0d,8'h18,8'h19,8'h1b,8'h11,8'h1f,8'h14,8'h20,8'h41,8'h2d,8'h3a,8'h4f,8'h7a,8'hc1,8'hea,8'hf8,8'hc4,8'h79,8'h6c,8'h63,8'h6c,8'h6f,8'h40,8'h67,8'hee,8'hfd,8'heb,8'h86,8'h2a,8'h26,8'h26,8'h26,8'h26,8'h25,8'h48,8'hce,8'hc6,8'h52,8'h63,8'h82,8'h66,8'h4e,8'h96,8'hfa,8'hed,8'h86,8'h2e,8'h25,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h47,8'h92,8'hdf,8'hf8,8'hff,8'hed,8'ha1,8'h66,8'h6f,8'h84,8'h84,8'h88,8'h70,8'h54,8'h4b,8'h6b,8'h9c,8'hc8,8'he7,8'hef,8'hf5,8'hff,8'hff,8'hd7,8'h63,8'h6e,8'h7c,8'h79,8'h7a,8'h81,8'h84,8'h80,8'h74,8'h4f,8'h49,8'h8c,8'he3,8'hff,8'hff,8'hf6,8'hd3,8'h82,8'h44,8'h26,8'h1f,8'h19,8'h1d,8'h19,8'h16,8'h14,8'h16,8'h1c,8'h1d,8'h0c,8'h12,8'h29,8'h2d,8'h3a,8'h29,8'h33,8'h36,8'h5a,8'h71,8'hab,8'h9f,8'h73,8'h78,8'h82,8'h88,8'h8d,8'hb4,8'hf1,8'hfa,8'h7e,8'h50,8'h74,8'h71,8'h72,8'h70,8'h6a,8'h6b,8'h4a,8'h3e,8'he3,8'hfb,8'h96,8'h23,8'h1a,8'h18,8'h1e,8'h23,8'h1b,8'h1c,8'h26,8'h2d,8'h2c,8'h2c,8'h11,8'h08,8'h11,8'h0d,8'h0f,8'h1a,8'h1a,8'h14,8'h15,8'h08,8'h11,8'h18,8'h14,8'h15,8'h07,8'h11,8'h11,8'h19,8'h18,8'h1b,8'h16,8'h24,8'h24,8'h2b,8'h27,8'h1f,8'h18,8'h21,8'h6c,8'hd9,8'hf8,8'hc4,8'h3c,8'h19,8'h15,8'h12,8'h19,8'h1b,8'h17,8'h14,8'h3c,8'h55,8'h1d,8'h16,8'h14,8'h1e,8'h1a,8'h11,8'h0f,8'h25,8'h49,8'h22,8'h1a,8'h0b,8'h10,8'h1d,8'h19,8'h1c,8'h12,8'h19,8'h14,8'h1b,8'h20,8'h17,8'h20,8'h17,8'h1f,8'h34,8'h66,8'hba,8'hee,8'hf2,8'hd6,8'h80,8'h49,8'h56,8'h46,8'h42,8'h97,8'hea,8'he6,8'h67,8'h28,8'h25,8'h26,8'h26,8'h25,8'h37,8'h9d,8'hda,8'h5f,8'h63,8'h8c,8'h6e,8'h40,8'h8d,8'hf2,8'hf7,8'h99,8'h33,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h28,8'h54,8'hbe,8'hf5,8'hff,8'hff,8'hd7,8'h77,8'h57,8'h73,8'h84,8'h89,8'h81,8'h5d,8'h4a,8'h6c,8'hac,8'heb,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfb,8'hfd,8'hb9,8'h5c,8'h6b,8'h75,8'h75,8'h79,8'h7d,8'h77,8'h64,8'h3c,8'h4e,8'hb3,8'hf4,8'hff,8'hfd,8'hec,8'had,8'h57,8'h26,8'h1f,8'h29,8'h24,8'h0c,8'h1f,8'h1b,8'h23,8'h22,8'h1f,8'h14,8'h0b,8'h12,8'h17,8'h20,8'h24,8'h21,8'h22,8'h44,8'h34,8'h44,8'h28,8'h4b,8'h37,8'h22,8'h24,8'h2a,8'h21,8'h23,8'h60,8'hec,8'hfd,8'h77,8'h4f,8'h7d,8'h73,8'h71,8'h71,8'h72,8'h6e,8'h4b,8'h43,8'he4,8'hf9,8'hb8,8'h4f,8'h25,8'h3c,8'h26,8'h26,8'h39,8'h20,8'h26,8'h25,8'h20,8'h2d,8'h1a,8'h1d,8'h16,8'h17,8'h11,8'h14,8'h0d,8'h0d,8'h0f,8'h0d,8'h12,8'h1b,8'h11,8'h14,8'h0c,8'h18,8'h0f,8'h16,8'h15,8'h13,8'h16,8'h34,8'h3a,8'h31,8'h26,8'h09,8'h23,8'h60,8'hd5,8'hfb,8'he1,8'h61,8'h0e,8'h14,8'h17,8'h10,8'h13,8'h14,8'h15,8'h1b,8'h35,8'h54,8'h20,8'h17,8'h15,8'h20,8'h1f,8'h1e,8'h21,8'h20,8'h23,8'h1e,8'h1a,8'h11,8'h11,8'h11,8'h12,8'h12,8'h14,8'h15,8'h15,8'h16,8'h0d,8'h14,8'h16,8'h19,8'h11,8'h19,8'h20,8'h3a,8'h7f,8'hce,8'hf9,8'hf0,8'had,8'h5d,8'h48,8'h47,8'h3b,8'h75,8'hda,8'hd7,8'h83,8'h3d,8'h26,8'h25,8'h2c,8'h83,8'he5,8'h88,8'h4c,8'h81,8'h7a,8'h42,8'h6d,8'heb,8'hff,8'hca,8'h49,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h00,8'h5b,8'hcb,8'hfb,8'hff,8'hfa,8'hb2,8'h5c,8'h64,8'h82,8'h83,8'h6e,8'h63,8'h4b,8'h66,8'hb9,8'hf5,8'hff,8'hff,8'hff,8'hf9,8'hee,8'he4,8'hec,8'hf8,8'hfa,8'h99,8'h5b,8'h70,8'h70,8'h77,8'h79,8'h78,8'h63,8'h4c,8'h74,8'hdb,8'hff,8'hfd,8'hf7,8'hd6,8'h7b,8'h2f,8'h1f,8'h16,8'h23,8'h26,8'h17,8'h10,8'h1b,8'h09,8'h27,8'h4b,8'h17,8'h10,8'h09,8'h1b,8'h1c,8'h20,8'h3f,8'h2a,8'h14,8'h26,8'h25,8'h2c,8'h14,8'h1b,8'h09,8'h40,8'h3a,8'h19,8'h1d,8'h24,8'h5a,8'hea,8'hfe,8'h71,8'h52,8'h7a,8'h75,8'h72,8'h76,8'h76,8'h73,8'h51,8'h46,8'he4,8'hf7,8'ha7,8'h38,8'h24,8'h2f,8'h2c,8'h26,8'h33,8'h27,8'h32,8'h2d,8'h20,8'h1f,8'h13,8'h23,8'h22,8'h13,8'h0a,8'h0f,8'h0c,8'h06,8'h0d,8'h12,8'h19,8'h19,8'h24,8'h4b,8'h45,8'h49,8'h1e,8'h17,8'h10,8'h0d,8'h1e,8'h1d,8'h18,8'h12,8'h0e,8'h12,8'h51,8'hce,8'hf9,8'hf0,8'h81,8'h20,8'h1a,8'h0b,8'h08,8'h11,8'h13,8'h14,8'h20,8'h28,8'h29,8'h3c,8'h14,8'h15,8'h14,8'h1b,8'h23,8'h41,8'h24,8'h16,8'h1e,8'h1e,8'h1d,8'h17,8'h14,8'h14,8'h15,8'h14,8'h10,8'h0c,8'h11,8'h13,8'h13,8'h10,8'h15,8'h19,8'h05,8'h09,8'h1a,8'h1c,8'h1c,8'h44,8'ha1,8'hec,8'hfc,8'hdc,8'h79,8'h46,8'h4c,8'h3a,8'h62,8'hcb,8'hea,8'had,8'h4e,8'h26,8'h58,8'hd8,8'hc2,8'h46,8'h74,8'h7f,8'h4f,8'h50,8'hd8,8'hff,8'hc8,8'h53,8'h28,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h29,8'h49,8'hbd,8'hfb,8'hff,8'hed,8'h8e,8'h50,8'h6e,8'h85,8'h82,8'h74,8'h56,8'h61,8'ha5,8'hef,8'hff,8'hff,8'hfb,8'hed,8'hcf,8'ha3,8'h75,8'h60,8'hba,8'hfd,8'hf2,8'h7a,8'h61,8'h78,8'h7b,8'h7d,8'h71,8'h4d,8'h48,8'ha0,8'hf5,8'hff,8'hfd,8'hed,8'hc2,8'h60,8'h23,8'h23,8'h23,8'h17,8'h18,8'h1f,8'h17,8'h1a,8'h18,8'h0d,8'h1e,8'h22,8'h0c,8'h1b,8'h14,8'h1a,8'h15,8'h29,8'h46,8'h1f,8'h20,8'h28,8'h24,8'h0f,8'h0e,8'h14,8'h12,8'h2d,8'h39,8'h1c,8'h2d,8'h4e,8'h65,8'hec,8'hfc,8'h6d,8'h58,8'h78,8'h73,8'h74,8'h79,8'h6f,8'h77,8'h5c,8'h48,8'he5,8'hfb,8'hbc,8'h2e,8'h15,8'h18,8'h2a,8'h2a,8'h29,8'h2d,8'h5c,8'h2b,8'h15,8'h23,8'h22,8'h2a,8'h26,8'h0b,8'h13,8'h16,8'h0a,8'h0a,8'h0f,8'h12,8'h14,8'h0c,8'h20,8'h6e,8'h6c,8'h31,8'h13,8'h0b,8'h15,8'h0e,8'h16,8'h14,8'h15,8'h0b,8'h0d,8'h47,8'hc4,8'hf8,8'hf7,8'hb3,8'h2c,8'h14,8'h20,8'h1b,8'h0c,8'h0c,8'h17,8'h15,8'h14,8'h22,8'h1e,8'h20,8'h1f,8'h1e,8'h19,8'h13,8'h0e,8'h16,8'h14,8'h19,8'h1d,8'h25,8'h24,8'h16,8'h10,8'h15,8'h18,8'h13,8'h12,8'h0f,8'h16,8'h15,8'h0f,8'h11,8'h0f,8'h17,8'h11,8'h06,8'h21,8'h3f,8'h1c,8'h14,8'h26,8'h65,8'hc4,8'hf8,8'hf3,8'ha3,8'h55,8'h43,8'h42,8'h4a,8'hae,8'hee,8'hbc,8'h62,8'hb7,8'he2,8'h60,8'h5f,8'h89,8'h5c,8'h42,8'hba,8'hff,8'he0,8'h67,8'h28,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h58,8'hc2,8'hf3,8'hff,8'he4,8'h7b,8'h5a,8'h73,8'h87,8'h83,8'h6a,8'h4f,8'h7b,8'hd7,8'hff,8'hff,8'hfd,8'he5,8'hbb,8'h7d,8'h47,8'h2c,8'h21,8'h36,8'hc3,8'hff,8'he3,8'h68,8'h6e,8'h81,8'h81,8'h65,8'h42,8'h54,8'hbc,8'hfe,8'hff,8'hfc,8'hdd,8'h88,8'h53,8'h3b,8'h24,8'h25,8'h22,8'h23,8'h21,8'h1d,8'h12,8'h12,8'h13,8'h10,8'h11,8'h1a,8'h15,8'h17,8'h19,8'h1b,8'h1e,8'h28,8'h2e,8'h0e,8'h24,8'h2c,8'h27,8'h32,8'h20,8'h1f,8'h1b,8'h2a,8'h46,8'h21,8'h24,8'h31,8'h6f,8'hf6,8'hfc,8'h6e,8'h5e,8'h77,8'h76,8'h76,8'h76,8'h72,8'h7b,8'h5b,8'h47,8'he6,8'hff,8'hb4,8'h25,8'h06,8'h14,8'h0e,8'h14,8'h12,8'h0f,8'h1c,8'h12,8'h15,8'h27,8'h39,8'h2c,8'h1e,8'h12,8'h24,8'h2c,8'h21,8'h0b,8'h14,8'h12,8'h0a,8'h05,8'h10,8'h4e,8'ha2,8'h3d,8'h1f,8'h12,8'h27,8'h2f,8'h1a,8'h15,8'h10,8'h0c,8'h41,8'hbe,8'hf5,8'hf9,8'hd0,8'h44,8'h14,8'h1c,8'h1a,8'h13,8'h0d,8'h10,8'h0d,8'h17,8'h1d,8'h22,8'h19,8'h0f,8'h15,8'h21,8'h1f,8'h1f,8'h17,8'h17,8'h23,8'h2a,8'h1c,8'h2f,8'h2b,8'h18,8'h19,8'h1a,8'h13,8'h11,8'h13,8'h17,8'h18,8'h0a,8'h0e,8'h0e,8'h11,8'h13,8'h1c,8'h25,8'h2c,8'h28,8'h28,8'h2d,8'h1f,8'h2c,8'h4a,8'h94,8'he4,8'hfa,8'hd0,8'h6d,8'h44,8'h40,8'h47,8'h8d,8'he4,8'hed,8'hf1,8'h8d,8'h47,8'h7e,8'h67,8'h3c,8'h96,8'hfa,8'hf4,8'h8e,8'h2c,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h29,8'h5b,8'hc6,8'hfc,8'hfb,8'hcd,8'h7f,8'h64,8'h7f,8'h86,8'h80,8'h60,8'h6d,8'ha4,8'hee,8'hff,8'hff,8'hdf,8'haa,8'h6e,8'h3c,8'h22,8'h1b,8'h20,8'h22,8'h52,8'hdd,8'hff,8'hc1,8'h60,8'h75,8'h73,8'h58,8'h58,8'h7f,8'hd6,8'hff,8'hff,8'he7,8'hab,8'h5b,8'h25,8'h45,8'h38,8'h25,8'h41,8'h24,8'h17,8'h26,8'h23,8'h21,8'h12,8'h1d,8'h16,8'h28,8'h3a,8'h1f,8'h20,8'h20,8'h3d,8'h40,8'h44,8'h23,8'h0b,8'h24,8'h2d,8'h2d,8'h4a,8'h22,8'h1f,8'h13,8'h13,8'h1e,8'h12,8'h14,8'h16,8'h72,8'hf7,8'hf9,8'h6e,8'h6a,8'h79,8'h79,8'h78,8'h78,8'h7b,8'h7c,8'h54,8'h49,8'he7,8'hff,8'had,8'h26,8'h14,8'h14,8'h09,8'h0f,8'h15,8'h14,8'h18,8'h17,8'h29,8'h3a,8'h34,8'h10,8'h25,8'h28,8'h2d,8'h21,8'h0f,8'h06,8'h0d,8'h12,8'h0a,8'h0c,8'h1b,8'h27,8'h96,8'hac,8'h3b,8'h0b,8'h3a,8'h6e,8'h22,8'h1a,8'h21,8'h51,8'hbc,8'hf6,8'hf8,8'hd5,8'h5a,8'h1d,8'h1e,8'h15,8'h14,8'h0a,8'h16,8'h14,8'h03,8'h22,8'h35,8'h23,8'h16,8'h16,8'h17,8'h19,8'h1d,8'h1d,8'h20,8'h27,8'h24,8'h30,8'h18,8'h1c,8'h17,8'h1f,8'h20,8'h19,8'h1e,8'h20,8'h1f,8'h20,8'h21,8'h32,8'h1b,8'h15,8'h0c,8'h2a,8'h29,8'h28,8'h2e,8'h0c,8'h2b,8'h34,8'h28,8'h37,8'h26,8'h2d,8'h65,8'hb6,8'heb,8'he7,8'h9f,8'h75,8'h42,8'h3b,8'h78,8'hb9,8'h92,8'h4b,8'h6c,8'h69,8'h49,8'h8a,8'hf3,8'hf5,8'hae,8'h45,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h42,8'hc0,8'hfd,8'hfd,8'hb7,8'h64,8'h6e,8'h86,8'h85,8'h7d,8'h4a,8'h65,8'hd6,8'hff,8'hfe,8'hf2,8'hc5,8'h65,8'h2a,8'h21,8'h1e,8'h20,8'h23,8'h20,8'h23,8'h73,8'hf1,8'hff,8'h94,8'h67,8'h77,8'h44,8'h51,8'hbb,8'hfd,8'hff,8'hf6,8'hd4,8'h74,8'h2c,8'h1b,8'h1f,8'h41,8'h2c,8'h20,8'h42,8'h37,8'h59,8'h74,8'h48,8'h46,8'h1c,8'h1a,8'h13,8'h2a,8'h3d,8'h21,8'h1c,8'h27,8'h63,8'hb8,8'hbb,8'h49,8'h1f,8'h18,8'h24,8'h27,8'h26,8'h14,8'h1b,8'h0f,8'h0e,8'h19,8'h1c,8'h16,8'h0f,8'h73,8'hf9,8'hf9,8'h6d,8'h68,8'h7c,8'h7f,8'h7e,8'h7f,8'h77,8'h72,8'h5b,8'h4b,8'hea,8'hfe,8'h96,8'h22,8'h1b,8'h18,8'h12,8'h0d,8'h0f,8'h14,8'h1f,8'h16,8'h27,8'h37,8'h26,8'h06,8'h27,8'h29,8'h12,8'h11,8'h0c,8'h0f,8'h0f,8'h12,8'h1f,8'h21,8'h13,8'h09,8'h4e,8'hd9,8'h9d,8'h1c,8'h3c,8'ha2,8'h37,8'h1c,8'h52,8'hcc,8'hf6,8'hfa,8'he6,8'h6c,8'h1f,8'h21,8'h10,8'h11,8'h22,8'h09,8'h16,8'h1a,8'h0e,8'h1c,8'h22,8'h19,8'h21,8'h20,8'h2c,8'h48,8'h25,8'h14,8'h1f,8'h26,8'h14,8'h1f,8'h1d,8'h18,8'h14,8'h20,8'h1f,8'h19,8'h20,8'h21,8'h1f,8'h22,8'h23,8'h33,8'h0b,8'h17,8'h16,8'h22,8'h20,8'h1d,8'h20,8'h0d,8'h1d,8'h1b,8'h1e,8'h23,8'h27,8'h31,8'h10,8'h53,8'h6f,8'hc9,8'hfa,8'he5,8'h7a,8'h3a,8'h42,8'h38,8'h30,8'h6a,8'h76,8'h44,8'h86,8'hf2,8'hf5,8'hae,8'h42,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3c,8'h95,8'hf4,8'hfc,8'hb2,8'h54,8'h6d,8'h86,8'h84,8'h76,8'h57,8'h64,8'hd8,8'hff,8'hfc,8'he6,8'h9c,8'h3f,8'h20,8'h1c,8'h1a,8'h1c,8'h2a,8'h33,8'h25,8'h28,8'h9c,8'hff,8'hf6,8'h71,8'h60,8'h48,8'h59,8'hcd,8'hff,8'hff,8'hf6,8'hc1,8'h5a,8'h25,8'h22,8'h23,8'h20,8'h2d,8'h2d,8'h36,8'h65,8'ha8,8'hd0,8'h88,8'h2a,8'h20,8'h1d,8'h15,8'h09,8'h24,8'h35,8'h1d,8'h23,8'h35,8'h71,8'he7,8'he5,8'h6d,8'h1b,8'h10,8'h1f,8'h23,8'h20,8'h1a,8'h17,8'h1f,8'h17,8'h14,8'h1a,8'h1b,8'h08,8'h70,8'hfa,8'hfb,8'h71,8'h64,8'h77,8'h79,8'h7e,8'h81,8'h79,8'h7d,8'h5b,8'h52,8'hee,8'hff,8'h94,8'h22,8'h19,8'h1d,8'h14,8'h0a,8'h0a,8'h10,8'h13,8'h1d,8'h19,8'h13,8'h21,8'h1b,8'h14,8'h11,8'h0f,8'h11,8'h28,8'h41,8'h26,8'h14,8'h35,8'h45,8'h13,8'h06,8'h25,8'ha4,8'he8,8'h65,8'h3a,8'hc0,8'h64,8'h4a,8'hc5,8'hf8,8'hf9,8'hf0,8'h8f,8'h25,8'h14,8'h1b,8'h0d,8'h18,8'h10,8'h09,8'h34,8'h2f,8'h11,8'h1a,8'h0a,8'h19,8'h21,8'h21,8'h3a,8'h5c,8'h25,8'h11,8'h10,8'h28,8'h2a,8'h22,8'h20,8'h16,8'h1f,8'h1f,8'h24,8'h36,8'h6a,8'h75,8'h30,8'h1f,8'h1a,8'h0c,8'h0b,8'h19,8'h19,8'h10,8'h13,8'h20,8'h21,8'h22,8'h1f,8'h1f,8'h25,8'h2f,8'h1c,8'h23,8'h0e,8'h1a,8'h25,8'h4b,8'ha9,8'hf4,8'hef,8'h93,8'h40,8'h52,8'h71,8'h7e,8'h49,8'h6c,8'heb,8'hfb,8'h9e,8'h3d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h54,8'hb5,8'hf3,8'hf7,8'ha3,8'h67,8'h7a,8'h8a,8'h85,8'h75,8'h54,8'h7d,8'hdf,8'hff,8'hfa,8'hcf,8'h77,8'h33,8'h21,8'h21,8'h22,8'h20,8'h21,8'h3b,8'h44,8'h2a,8'h3d,8'hc6,8'hff,8'hdc,8'h40,8'h47,8'h8a,8'hdf,8'hff,8'hfe,8'hdf,8'hb7,8'h4d,8'h23,8'h21,8'h23,8'h22,8'h2f,8'h60,8'h93,8'hbc,8'he3,8'hf4,8'hb0,8'h53,8'h23,8'h10,8'h1a,8'h0f,8'h0f,8'h22,8'h20,8'h10,8'h21,8'h18,8'h39,8'h92,8'h9f,8'h41,8'h14,8'h17,8'h15,8'h1b,8'h1f,8'h1c,8'h14,8'h13,8'h1f,8'h23,8'h1a,8'h0f,8'h09,8'h74,8'hfb,8'hfa,8'h6f,8'h65,8'h79,8'h79,8'h7c,8'h79,8'h74,8'h7e,8'h5d,8'h58,8'hf2,8'hff,8'ha5,8'h2b,8'h25,8'h1f,8'h1a,8'h1b,8'h19,8'h20,8'h09,8'h13,8'h12,8'h0b,8'h19,8'h22,8'h1a,8'h11,8'h0c,8'h05,8'h27,8'h4b,8'h23,8'h14,8'h22,8'h22,8'h09,8'h11,8'h18,8'h5a,8'hdf,8'hd2,8'h9e,8'hde,8'hca,8'hcb,8'hf5,8'hf7,8'hf3,8'h9d,8'h2d,8'h12,8'h14,8'h18,8'h14,8'h17,8'h0e,8'h1a,8'h29,8'h21,8'h10,8'h22,8'h19,8'h16,8'h26,8'h26,8'h28,8'h22,8'h22,8'h27,8'h1f,8'h27,8'h21,8'h1f,8'h1c,8'h20,8'h33,8'h62,8'h93,8'hc5,8'hed,8'hcf,8'h4f,8'h17,8'h17,8'h13,8'h11,8'h14,8'h12,8'h0e,8'h13,8'h17,8'h24,8'h38,8'h1d,8'h18,8'h10,8'h1d,8'h0f,8'h14,8'h1b,8'h26,8'h39,8'h2d,8'h45,8'hd7,8'hff,8'hd7,8'h4b,8'h6c,8'h83,8'h50,8'h7c,8'he1,8'hfd,8'hba,8'h42,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h4a,8'hc5,8'hff,8'hf9,8'ha3,8'h4c,8'h80,8'h8f,8'h86,8'h83,8'h58,8'h6b,8'he4,8'hff,8'hfc,8'hd4,8'h66,8'h26,8'h1b,8'h1f,8'h20,8'h21,8'h22,8'h20,8'h29,8'h34,8'h32,8'h54,8'he6,8'hff,8'ha6,8'h43,8'hab,8'hfc,8'hff,8'hfa,8'hd0,8'h67,8'h30,8'h20,8'h22,8'h22,8'h30,8'h56,8'ha0,8'hd9,8'hf6,8'hfe,8'hff,8'hdd,8'h58,8'h23,8'h18,8'h17,8'h19,8'h18,8'h17,8'h1a,8'h0f,8'h10,8'h1e,8'h08,8'h0f,8'h32,8'h3d,8'h29,8'h21,8'h14,8'h17,8'h1a,8'h1c,8'h1f,8'h0a,8'h01,8'h22,8'h40,8'h20,8'h27,8'h2f,8'h79,8'hfc,8'hf9,8'h6d,8'h67,8'h77,8'h7b,8'h7a,8'h7b,8'h77,8'h7b,8'h5b,8'h61,8'hf5,8'hff,8'h98,8'h36,8'h40,8'h26,8'h10,8'h1b,8'h10,8'h13,8'h0c,8'h0d,8'h0b,8'h08,8'h09,8'h10,8'h27,8'h24,8'h0f,8'h0b,8'h1d,8'h51,8'h2c,8'h1d,8'h17,8'h14,8'h1c,8'h16,8'h0b,8'h24,8'h9f,8'hf6,8'hf6,8'hf5,8'hf8,8'hf9,8'hf7,8'hf8,8'hcb,8'h37,8'h25,8'h37,8'h4e,8'h47,8'h1d,8'h10,8'h1a,8'h14,8'h0d,8'h05,8'h0e,8'h13,8'h1e,8'h11,8'h21,8'h25,8'h20,8'h18,8'h1f,8'h24,8'h24,8'h20,8'h10,8'h24,8'h3b,8'h6f,8'hb0,8'he5,8'hf9,8'hff,8'hec,8'h7a,8'h25,8'h1b,8'h14,8'h14,8'h0e,8'h0f,8'h14,8'h19,8'h2e,8'h22,8'h23,8'h4c,8'h14,8'h0e,8'h13,8'h1a,8'h15,8'h1d,8'h1f,8'h1f,8'h22,8'h21,8'h7b,8'hf4,8'hf5,8'h78,8'h4b,8'h7d,8'h48,8'h63,8'he8,8'hff,8'hc8,8'h4f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h34,8'ha2,8'hf9,8'hfd,8'hbe,8'h5a,8'h6f,8'h86,8'h83,8'h85,8'h6a,8'h5d,8'hcf,8'hff,8'hff,8'hde,8'h6b,8'h29,8'h22,8'h1f,8'h1b,8'h20,8'h22,8'h24,8'h24,8'h20,8'h21,8'h23,8'h77,8'hf6,8'hff,8'h9c,8'hb1,8'hff,8'hff,8'hf3,8'hc9,8'h61,8'h20,8'h0f,8'h27,8'h37,8'h5e,8'ha3,8'hd9,8'hf4,8'hfe,8'hff,8'hfe,8'hf4,8'h91,8'h37,8'h44,8'h1b,8'h1d,8'h1f,8'h1f,8'h1b,8'h18,8'h14,8'h17,8'h15,8'h07,8'h01,8'h14,8'h22,8'h10,8'h16,8'h19,8'h18,8'h1f,8'h1f,8'h1f,8'h18,8'h12,8'h22,8'h28,8'h20,8'h27,8'h2b,8'h78,8'hfd,8'hf4,8'h6a,8'h66,8'h75,8'h78,8'h7a,8'h7e,8'h82,8'h7b,8'h5b,8'h63,8'hf6,8'hfa,8'h90,8'h25,8'h22,8'h1d,8'h25,8'h2a,8'h19,8'h20,8'h21,8'h14,8'h0e,8'h03,8'h0a,8'h16,8'h3e,8'h42,8'h11,8'h18,8'h15,8'h22,8'h04,8'h07,8'h0e,8'h19,8'h1a,8'h1b,8'h0c,8'h17,8'h61,8'he6,8'hf8,8'hf7,8'hf7,8'hf7,8'hf7,8'hf7,8'hcc,8'h8a,8'h9c,8'h9b,8'h67,8'h2e,8'h19,8'h19,8'h17,8'h0b,8'h10,8'h1f,8'h24,8'h21,8'h1b,8'h1f,8'h21,8'h24,8'h1a,8'h15,8'h1e,8'h2a,8'h41,8'h32,8'h46,8'h83,8'hc4,8'hea,8'hfc,8'hff,8'hff,8'hf2,8'h9d,8'h2d,8'h19,8'h1a,8'h10,8'h0e,8'h0a,8'h14,8'h1b,8'h19,8'h29,8'h20,8'h23,8'h29,8'h16,8'h18,8'h21,8'h21,8'h15,8'h12,8'h1b,8'h12,8'h1f,8'h5c,8'hdf,8'hff,8'ha6,8'h3d,8'h64,8'h51,8'h5f,8'hd8,8'hff,8'hde,8'h66,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2a,8'h79,8'hec,8'hfd,8'hb1,8'h64,8'h85,8'h8c,8'h85,8'h82,8'h71,8'h62,8'hc4,8'hff,8'hfb,8'hdd,8'h6e,8'h23,8'h22,8'h23,8'h20,8'h20,8'h22,8'h30,8'h36,8'h45,8'h29,8'h24,8'h29,8'haf,8'hff,8'hff,8'hf6,8'hfd,8'hfd,8'hf1,8'hb6,8'h4d,8'h24,8'h27,8'h4a,8'h8e,8'hc5,8'he5,8'hf9,8'hff,8'hff,8'hff,8'hff,8'hf9,8'hbb,8'h3e,8'h20,8'h28,8'h1f,8'h1f,8'h20,8'h20,8'h1b,8'h15,8'h16,8'h16,8'h1c,8'h20,8'h25,8'h3f,8'h51,8'h34,8'h29,8'h21,8'h27,8'h4b,8'h2e,8'h34,8'h37,8'h33,8'h30,8'h29,8'h20,8'h1d,8'h15,8'h7b,8'hff,8'hf1,8'h65,8'h6c,8'h7a,8'h7a,8'h7b,8'h7a,8'h7d,8'h7b,8'h59,8'h64,8'hf6,8'hf7,8'h8f,8'h27,8'h30,8'h35,8'h2f,8'h33,8'h2b,8'h2b,8'h44,8'h22,8'h13,8'h13,8'h1b,8'h1e,8'h14,8'h0d,8'h04,8'h0c,8'h23,8'h39,8'h4a,8'h63,8'h76,8'h7e,8'h81,8'h83,8'h83,8'h93,8'hc3,8'hf0,8'hf7,8'hf7,8'hf7,8'hf7,8'hf7,8'hf7,8'hf0,8'ha5,8'h52,8'h2e,8'h10,8'h0e,8'h1b,8'h14,8'h0d,8'h12,8'h22,8'h23,8'h43,8'h31,8'h1d,8'h1f,8'h20,8'h24,8'h21,8'h2a,8'h43,8'h73,8'hab,8'hc8,8'he0,8'hf4,8'hfa,8'hff,8'hff,8'hff,8'hf5,8'ha4,8'h3b,8'h1d,8'h23,8'h15,8'h10,8'h11,8'h15,8'h24,8'h26,8'h1f,8'h0b,8'h03,8'h36,8'h3d,8'h2d,8'h0b,8'h2f,8'h27,8'h1f,8'h1f,8'h20,8'h16,8'h56,8'hd5,8'hff,8'hb7,8'h4a,8'h5f,8'h44,8'h61,8'hd8,8'hff,8'hd9,8'h64,8'h2a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h28,8'h66,8'hda,8'hff,8'hd8,8'h63,8'h76,8'h8e,8'h80,8'h85,8'h75,8'h52,8'h92,8'hfe,8'hff,8'he9,8'h88,8'h26,8'h16,8'h23,8'h22,8'h1f,8'h17,8'h22,8'h24,8'h31,8'h42,8'h40,8'h26,8'h3a,8'hd3,8'hff,8'hff,8'hff,8'hff,8'hea,8'h9e,8'h4d,8'h25,8'h4b,8'h94,8'hd6,8'hf4,8'hfe,8'hff,8'hff,8'hf1,8'hff,8'hff,8'hff,8'he5,8'h63,8'h14,8'h22,8'h26,8'h21,8'h20,8'h1f,8'h20,8'h14,8'h0b,8'h19,8'h26,8'h43,8'h6f,8'h98,8'hbe,8'hcb,8'hbe,8'had,8'h85,8'h66,8'h58,8'h2f,8'h4b,8'h34,8'h28,8'h1c,8'h16,8'h10,8'h0d,8'h0f,8'h85,8'hff,8'he4,8'h56,8'h6a,8'h7d,8'h7d,8'h7b,8'h79,8'h82,8'h81,8'h5b,8'h6a,8'hf9,8'hf9,8'ha5,8'h43,8'h25,8'h3a,8'h33,8'h36,8'h39,8'h27,8'h20,8'h17,8'h12,8'h1a,8'h20,8'h16,8'h07,8'h11,8'h27,8'h27,8'h2a,8'h40,8'h52,8'h73,8'h90,8'ha8,8'hc2,8'hd2,8'he0,8'hed,8'hf7,8'hf7,8'hf7,8'hf7,8'hf7,8'hf7,8'hf8,8'hf9,8'hf4,8'h8d,8'h45,8'h44,8'h3a,8'h30,8'h26,8'h1d,8'h18,8'h19,8'h17,8'h1f,8'h1f,8'h14,8'h18,8'h1f,8'h25,8'h42,8'h74,8'ha6,8'hd0,8'hef,8'hfc,8'hff,8'hf0,8'hc0,8'h9e,8'hec,8'hff,8'hfc,8'hc1,8'h42,8'h14,8'h17,8'h1e,8'h0e,8'h13,8'h14,8'h09,8'h20,8'h45,8'h26,8'h11,8'h15,8'h22,8'h25,8'h22,8'h10,8'h40,8'h2d,8'h1a,8'h1b,8'h27,8'h4c,8'hc1,8'hff,8'hdf,8'h4f,8'h51,8'h48,8'h4c,8'hcd,8'hff,8'hee,8'h73,8'h29,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h49,8'hca,8'hff,8'he7,8'h85,8'h6b,8'h88,8'h84,8'h82,8'h80,8'h69,8'h6a,8'he2,8'hff,8'hf3,8'hb1,8'h41,8'h20,8'h21,8'h22,8'h21,8'h1f,8'h1d,8'h26,8'h36,8'h3a,8'h2e,8'h25,8'h1f,8'h5d,8'hea,8'hff,8'hff,8'hfc,8'hd8,8'h96,8'h58,8'h5d,8'h91,8'hd6,8'hf9,8'hff,8'hfa,8'he1,8'hc4,8'h8b,8'h90,8'hf6,8'hff,8'hf6,8'hb5,8'h30,8'h23,8'h2e,8'h2d,8'h18,8'h20,8'h14,8'h21,8'h37,8'h4c,8'h6b,8'h9d,8'hce,8'heb,8'hf8,8'hff,8'hff,8'hff,8'hff,8'hf4,8'hd9,8'h9b,8'h5d,8'h31,8'h10,8'h14,8'h1f,8'h1c,8'h1c,8'h32,8'h32,8'h91,8'hff,8'hda,8'h57,8'h7a,8'h7a,8'h7d,8'h7c,8'h79,8'h7b,8'h79,8'h5f,8'h67,8'hf6,8'hfd,8'haa,8'h47,8'h33,8'h35,8'h2d,8'h41,8'h31,8'h2a,8'h1f,8'h19,8'h0b,8'h21,8'h36,8'h48,8'h5e,8'h85,8'hb9,8'hb8,8'h94,8'h71,8'h5b,8'h54,8'h5b,8'h5b,8'h4b,8'h3f,8'h62,8'hba,8'hf2,8'hf8,8'hf7,8'hf7,8'hf7,8'hf7,8'heb,8'hd0,8'hc2,8'hac,8'h98,8'h91,8'h84,8'h72,8'h45,8'h23,8'h12,8'h11,8'h0a,8'h1e,8'h2f,8'h48,8'h59,8'h75,8'ha4,8'hd2,8'hef,8'hff,8'hff,8'he7,8'hce,8'hba,8'h75,8'h3e,8'h85,8'hf2,8'hff,8'hdb,8'h5e,8'h1d,8'h17,8'h25,8'h2b,8'h23,8'h11,8'h0c,8'h0f,8'h14,8'h29,8'h29,8'h1f,8'h24,8'h27,8'h10,8'h12,8'h1d,8'h29,8'h5a,8'h68,8'h69,8'h98,8'hd1,8'hfa,8'he9,8'h73,8'h3f,8'h4f,8'h4a,8'hbd,8'hff,8'hff,8'hef,8'h8c,8'h38,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h34,8'ha6,8'hfc,8'hf2,8'h82,8'h6f,8'h88,8'h82,8'h85,8'h84,8'h77,8'h5b,8'hc1,8'hff,8'hff,8'hd3,8'h51,8'h20,8'h23,8'h23,8'h22,8'h21,8'h20,8'h1f,8'h21,8'h26,8'h26,8'h28,8'h21,8'h23,8'h93,8'hfc,8'hff,8'hfe,8'hd2,8'h7d,8'h88,8'hc8,8'he6,8'hf5,8'hff,8'hfe,8'hdc,8'h8c,8'h4a,8'h32,8'h2c,8'hb4,8'hff,8'hff,8'hcf,8'h6f,8'h42,8'h2d,8'h27,8'h21,8'h20,8'h33,8'h55,8'h8e,8'hca,8'he2,8'hed,8'hfb,8'hff,8'hfd,8'hf6,8'hec,8'he7,8'he7,8'hf7,8'hff,8'hff,8'hf7,8'he1,8'h8c,8'h2d,8'h12,8'h20,8'h1c,8'h22,8'h40,8'h31,8'h96,8'hff,8'hd4,8'h55,8'h7e,8'h79,8'h78,8'h77,8'h77,8'h7e,8'h7d,8'h60,8'h66,8'hf6,8'hff,8'h8e,8'h37,8'h31,8'h27,8'h3b,8'h4e,8'h40,8'h20,8'h27,8'h32,8'h57,8'h8d,8'hc1,8'hdf,8'hed,8'hf8,8'hff,8'hfb,8'he0,8'hae,8'h85,8'h73,8'h72,8'h60,8'h2f,8'h40,8'h80,8'hb9,8'hec,8'hf8,8'hf7,8'hf7,8'hf8,8'hf5,8'h9d,8'h35,8'h29,8'h27,8'h2b,8'h32,8'h3f,8'h45,8'h25,8'h20,8'h21,8'h33,8'h4f,8'h77,8'hb8,8'hde,8'hea,8'hf3,8'hfc,8'hfe,8'hed,8'hcd,8'h97,8'h61,8'h55,8'h5b,8'h35,8'h72,8'hed,8'hfe,8'hfd,8'hc6,8'h3e,8'h20,8'h1e,8'h23,8'h34,8'h2e,8'h0e,8'h12,8'h22,8'h28,8'h24,8'h42,8'h27,8'h3a,8'h32,8'h23,8'h36,8'h55,8'h85,8'hca,8'he6,8'hef,8'hfb,8'hff,8'hef,8'h75,8'h3d,8'h40,8'h1d,8'h46,8'h99,8'hd6,8'hfb,8'hff,8'hf1,8'haf,8'h47,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h28,8'h72,8'hea,8'hff,8'hac,8'h55,8'h83,8'h8f,8'h8b,8'h83,8'h86,8'h65,8'h74,8'hf7,8'hff,8'hee,8'h84,8'h22,8'h1c,8'h23,8'h23,8'h21,8'h21,8'h20,8'h22,8'h2a,8'h24,8'h21,8'h23,8'h20,8'h30,8'hc6,8'hff,8'hfe,8'hf5,8'hc7,8'hc6,8'hec,8'hfb,8'hfd,8'hf5,8'hd5,8'h85,8'h47,8'h48,8'h63,8'h45,8'h69,8'hf5,8'hff,8'hef,8'h87,8'h2f,8'h41,8'h2a,8'h34,8'h50,8'h81,8'hbd,8'he6,8'hfa,8'hfd,8'hfe,8'hf8,8'he1,8'hba,8'h87,8'h68,8'h4e,8'h46,8'h4a,8'h65,8'ha2,8'he9,8'hff,8'hff,8'hea,8'h87,8'h22,8'h0d,8'h15,8'h0f,8'h17,8'h22,8'h9a,8'hff,8'hd4,8'h56,8'h7a,8'h77,8'h79,8'h77,8'h7e,8'h7f,8'h83,8'h66,8'h65,8'hf7,8'hff,8'h97,8'h53,8'h2b,8'h22,8'h2f,8'h50,8'h6d,8'h66,8'h92,8'hc2,8'he7,8'hfa,8'hff,8'hff,8'hfc,8'he7,8'hb6,8'h76,8'h4a,8'h38,8'h36,8'h37,8'h26,8'h25,8'h27,8'h36,8'h2b,8'h43,8'hc9,8'hfa,8'hf9,8'hf7,8'hf8,8'hf5,8'h8b,8'h16,8'h0c,8'h11,8'h19,8'h15,8'h30,8'h4e,8'h3c,8'h66,8'h97,8'hc8,8'he5,8'hf5,8'hfb,8'hfc,8'hf9,8'he9,8'hc9,8'h9c,8'h65,8'h48,8'h49,8'h57,8'h62,8'h49,8'h61,8'he2,8'hff,8'hff,8'hfc,8'hf0,8'h90,8'h27,8'h17,8'h13,8'h10,8'h1b,8'h20,8'h1b,8'h26,8'h3b,8'h25,8'h22,8'h23,8'h35,8'h55,8'h7b,8'hbc,8'he2,8'hf2,8'hfd,8'hff,8'hff,8'hf4,8'hd1,8'h7a,8'h32,8'h4b,8'h31,8'h2d,8'h34,8'h36,8'h41,8'h86,8'he6,8'hff,8'hf7,8'haa,8'h3c,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h4f,8'hcd,8'hff,8'hcc,8'h62,8'h74,8'h8c,8'h89,8'h87,8'h88,8'h7a,8'h58,8'hba,8'hff,8'hfd,8'hbc,8'h40,8'h21,8'h20,8'h20,8'h21,8'h20,8'h22,8'h20,8'h23,8'h23,8'h21,8'h22,8'h23,8'h1d,8'h52,8'he3,8'hff,8'hfe,8'hf9,8'hf4,8'hf9,8'hf9,8'hdc,8'ha5,8'h80,8'h58,8'h48,8'h5f,8'h81,8'h67,8'h50,8'hc8,8'hff,8'hf9,8'hae,8'h56,8'h57,8'h78,8'h8a,8'hb9,8'hdd,8'hf4,8'hff,8'hff,8'he1,8'hb2,8'h95,8'h82,8'h60,8'h4b,8'h43,8'h42,8'h44,8'h4d,8'h4f,8'h43,8'h4b,8'h72,8'hb8,8'hf8,8'hff,8'he3,8'h6e,8'h18,8'h09,8'h11,8'h1c,8'h25,8'ha9,8'hff,8'hd5,8'h5c,8'h7d,8'h7a,8'h7d,8'h7e,8'h82,8'h81,8'h86,8'h6b,8'h63,8'hf4,8'hff,8'ha2,8'h41,8'h5c,8'h78,8'h86,8'ha5,8'hce,8'heb,8'hfd,8'hff,8'hfa,8'he0,8'hb2,8'h97,8'h87,8'h68,8'h50,8'h40,8'h4c,8'h66,8'h6f,8'h6e,8'h64,8'h68,8'h6a,8'h55,8'h26,8'h65,8'he4,8'he6,8'hbe,8'hdd,8'hc3,8'he9,8'hb1,8'h2d,8'h25,8'h22,8'h23,8'h49,8'h84,8'h9e,8'hc2,8'he8,8'hf9,8'hff,8'hfa,8'he4,8'hb8,8'h98,8'h94,8'h74,8'h5d,8'h4e,8'h51,8'h66,8'h70,8'h67,8'h51,8'h62,8'hcb,8'hf5,8'he5,8'he8,8'hfb,8'hfe,8'hc4,8'h36,8'h15,8'h1c,8'h18,8'h29,8'h37,8'h1c,8'h30,8'h2a,8'h46,8'h70,8'h88,8'hab,8'hd8,8'hef,8'hfc,8'hff,8'hfa,8'hdf,8'hb6,8'h98,8'h75,8'h50,8'h48,8'h55,8'h61,8'h61,8'h72,8'h74,8'h73,8'h60,8'h43,8'h67,8'hd8,8'hff,8'hec,8'h86,8'h2d,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3a,8'hab,8'hfa,8'hf2,8'h71,8'h67,8'h91,8'h85,8'h83,8'h85,8'h8d,8'h68,8'h6c,8'hf3,8'hff,8'he5,8'h6d,8'h21,8'h23,8'h21,8'h20,8'h22,8'h22,8'h20,8'h1f,8'h20,8'h20,8'h21,8'h22,8'h23,8'h3d,8'h9e,8'hf8,8'hff,8'hfd,8'hff,8'hff,8'he2,8'h96,8'h50,8'h3c,8'h55,8'h6a,8'h81,8'h8d,8'h7f,8'h45,8'h9b,8'hff,8'hfd,8'hf1,8'hb9,8'hb0,8'hdf,8'hf4,8'hfc,8'hff,8'hff,8'hf0,8'hc9,8'h8d,8'h58,8'h43,8'h47,8'h59,8'h66,8'h6e,8'h77,8'h73,8'h75,8'h7c,8'h77,8'h72,8'h6e,8'h5d,8'h49,8'had,8'hff,8'hff,8'hca,8'h3f,8'h0b,8'h1b,8'h14,8'h21,8'hb0,8'hff,8'hd4,8'h5e,8'h79,8'h7d,8'h83,8'h83,8'h83,8'h85,8'h8a,8'h6a,8'h67,8'hf4,8'hff,8'hd7,8'hb8,8'hde,8'hf0,8'hfb,8'hff,8'hff,8'hff,8'he6,8'hb4,8'h77,8'h4b,8'h3b,8'h47,8'h57,8'h60,8'h6a,8'h6a,8'h69,8'h72,8'h73,8'h76,8'h7b,8'h7f,8'h79,8'h5b,8'h63,8'hd5,8'he0,8'h6c,8'h5b,8'hc2,8'h62,8'hb6,8'hc0,8'h3d,8'h39,8'h23,8'h5f,8'hc9,8'hf2,8'hfc,8'hff,8'hfe,8'hef,8'hc1,8'h82,8'h5a,8'h4a,8'h4a,8'h56,8'h5c,8'h65,8'h6c,8'h6b,8'h6e,8'h71,8'h6c,8'h3a,8'h58,8'h84,8'h62,8'h4c,8'h54,8'hc7,8'hff,8'hce,8'h41,8'h1c,8'h1e,8'h17,8'h24,8'h2f,8'h3a,8'h75,8'h9f,8'hd0,8'hed,8'hfa,8'hfb,8'hff,8'hff,8'hf9,8'hd0,8'h8b,8'h50,8'h3a,8'h43,8'h54,8'h5d,8'h6b,8'h6a,8'h69,8'h6b,8'h76,8'h7b,8'h7d,8'h85,8'h80,8'h4a,8'h6b,8'hf0,8'hff,8'hd0,8'h45,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h29,8'h78,8'hed,8'hff,8'hb3,8'h55,8'h81,8'h8b,8'h81,8'h85,8'h7f,8'h7f,8'h56,8'ha8,8'hff,8'hff,8'hbe,8'h39,8'h21,8'h26,8'h21,8'h21,8'h22,8'h23,8'h36,8'h29,8'h21,8'h23,8'h23,8'h2d,8'h63,8'hb0,8'hee,8'hff,8'hfe,8'hff,8'hfd,8'ha7,8'h4e,8'h45,8'h53,8'h74,8'h83,8'h83,8'h83,8'h81,8'h59,8'h63,8'hea,8'hff,8'hf6,8'hf5,8'hf1,8'hf9,8'hf5,8'hf4,8'hec,8'hc7,8'h92,8'h62,8'h47,8'h48,8'h57,8'h69,8'h6e,8'h70,8'h70,8'h71,8'h73,8'h76,8'h74,8'h7d,8'h78,8'h75,8'h77,8'h74,8'h43,8'h50,8'he7,8'hff,8'he9,8'h5b,8'h17,8'h1d,8'h0f,8'h26,8'hb6,8'hff,8'hd0,8'h61,8'h78,8'h77,8'h7f,8'h84,8'h89,8'h85,8'h8b,8'h6c,8'h6a,8'hf3,8'hfd,8'hfb,8'hfd,8'hfd,8'hf9,8'hfa,8'hea,8'hc0,8'h86,8'h4e,8'h3c,8'h42,8'h58,8'h68,8'h71,8'h6e,8'h70,8'h6c,8'h6a,8'h6c,8'h71,8'h74,8'h74,8'h74,8'h7a,8'h6c,8'h54,8'hae,8'hd1,8'h7c,8'h5d,8'hb1,8'hda,8'h43,8'h6d,8'hb6,8'h31,8'h17,8'h4c,8'hd3,8'hfc,8'hfb,8'hf7,8'he5,8'hab,8'h66,8'h40,8'h3b,8'h4f,8'h63,8'h62,8'h64,8'h63,8'h66,8'h67,8'h65,8'h71,8'h75,8'h76,8'h4e,8'h2f,8'h3e,8'h47,8'h46,8'h36,8'h97,8'hff,8'hcd,8'h41,8'h20,8'h24,8'h34,8'h58,8'h8a,8'hc3,8'he5,8'hf7,8'hff,8'hfd,8'hfb,8'hf7,8'he4,8'hb5,8'h6e,8'h44,8'h3f,8'h4f,8'h61,8'h69,8'h6e,8'h6c,8'h68,8'h66,8'h64,8'h65,8'h6d,8'h74,8'h79,8'h7f,8'h88,8'h70,8'h40,8'hba,8'hff,8'hea,8'h61,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h4d,8'hd0,8'hff,8'hd4,8'h66,8'h73,8'h83,8'h82,8'h87,8'h81,8'h7d,8'h69,8'h60,8'he1,8'hff,8'hf2,8'h7e,8'h22,8'h21,8'h20,8'h1f,8'h30,8'h43,8'h21,8'h2c,8'h23,8'h15,8'h22,8'h22,8'h32,8'h66,8'h84,8'hc0,8'he6,8'hfc,8'hff,8'hfb,8'h93,8'h35,8'h6c,8'h77,8'h81,8'h7f,8'h81,8'h87,8'h6a,8'h48,8'hbe,8'hff,8'hfb,8'hfc,8'hf9,8'he1,8'hb9,8'h7c,8'h5d,8'h5a,8'h51,8'h55,8'h59,8'h6c,8'h7f,8'h72,8'h6d,8'h70,8'h6b,8'h6a,8'h6b,8'h6b,8'h6e,8'h73,8'h77,8'h79,8'h79,8'h77,8'h73,8'h6b,8'h4c,8'hae,8'hff,8'hf6,8'h71,8'h2c,8'h24,8'h3b,8'h33,8'hb8,8'hff,8'hcd,8'h58,8'h72,8'h79,8'h7f,8'h85,8'h87,8'h8a,8'h92,8'h6d,8'h72,8'hfa,8'hff,8'hff,8'hea,8'hb5,8'h76,8'h56,8'h40,8'h32,8'h4a,8'h51,8'h65,8'h78,8'h7a,8'h72,8'h6d,8'h6e,8'h72,8'h6d,8'h6e,8'h6e,8'h6e,8'h6e,8'h73,8'h79,8'h71,8'h4d,8'h84,8'h95,8'h48,8'h73,8'he0,8'hf9,8'hce,8'h2f,8'h2d,8'h8c,8'h45,8'h23,8'haa,8'hfd,8'hff,8'hc0,8'h70,8'h5f,8'h56,8'h58,8'h66,8'h6c,8'h6c,8'h6b,8'h67,8'h6a,8'h6a,8'h6d,8'h70,8'h70,8'h73,8'h75,8'h79,8'h74,8'h6c,8'h6d,8'h72,8'h6a,8'h4a,8'ha4,8'hff,8'hc8,8'h3e,8'h58,8'ha8,8'hc6,8'he2,8'hf6,8'hfa,8'hfe,8'hff,8'he4,8'hb4,8'h76,8'h5e,8'h57,8'h52,8'h53,8'h5b,8'h67,8'h6f,8'h6c,8'h67,8'h6e,8'h6b,8'h68,8'h68,8'h68,8'h6a,8'h6c,8'h73,8'h75,8'h77,8'h82,8'h84,8'h44,8'h82,8'hfe,8'hfa,8'h81,8'h29,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h32,8'ha2,8'hfb,8'hf9,8'h88,8'h63,8'h81,8'h7d,8'h7f,8'h81,8'h7a,8'h7a,8'h5f,8'h82,8'hfd,8'hff,8'hd5,8'h4e,8'h1f,8'h21,8'h27,8'h28,8'h32,8'h4f,8'h36,8'h22,8'h20,8'h19,8'h1a,8'h24,8'h25,8'h25,8'h2a,8'h37,8'h5f,8'hc0,8'hf7,8'hff,8'hf0,8'h74,8'h61,8'h77,8'h80,8'h7d,8'h7d,8'h80,8'h46,8'h78,8'hfd,8'hff,8'hff,8'hff,8'he1,8'h83,8'h4a,8'h34,8'h2d,8'h44,8'h57,8'h56,8'h4f,8'h50,8'h61,8'h74,8'h6e,8'h72,8'h73,8'h6e,8'h6f,8'h6e,8'h6c,8'h70,8'h71,8'h75,8'h7f,8'h77,8'h77,8'h7a,8'h53,8'h86,8'hff,8'hf9,8'h7c,8'h40,8'h28,8'h46,8'h3a,8'hbc,8'hff,8'hcc,8'h5a,8'h7c,8'h80,8'h81,8'h87,8'h87,8'h86,8'h8e,8'h69,8'h76,8'hff,8'hff,8'hff,8'hcd,8'h80,8'h5e,8'h4d,8'h45,8'h43,8'h43,8'h3d,8'h37,8'h3a,8'h53,8'h7f,8'h74,8'h70,8'h74,8'h72,8'h6d,8'h6d,8'h72,8'h6e,8'h74,8'h72,8'h4d,8'h51,8'h76,8'h48,8'h3c,8'h9b,8'hfc,8'hf6,8'h90,8'h23,8'h1b,8'h4c,8'h40,8'h43,8'hde,8'hff,8'hd0,8'h42,8'h40,8'h66,8'h75,8'h71,8'h6e,8'h6d,8'h6e,8'h6a,8'h68,8'h71,8'h71,8'h70,8'h6e,8'h71,8'h73,8'h73,8'h76,8'h6e,8'h70,8'h6e,8'h6f,8'h6b,8'h46,8'hb1,8'hff,8'hbd,8'h44,8'had,8'hfe,8'hff,8'hfc,8'hff,8'hff,8'hff,8'hf9,8'ha5,8'h5f,8'h41,8'h36,8'h43,8'h4a,8'h49,8'h4c,8'h59,8'h69,8'h66,8'h6a,8'h6e,8'h6a,8'h6e,8'h6c,8'h6c,8'h6c,8'h6a,8'h6d,8'h73,8'h7b,8'h81,8'h87,8'h4e,8'h6b,8'hf7,8'hff,8'h89,8'h2a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h5d,8'he1,8'hff,8'hcc,8'h60,8'h77,8'h84,8'h7f,8'h80,8'h7f,8'h80,8'h78,8'h54,8'had,8'hff,8'hfc,8'haa,8'h31,8'h1f,8'h20,8'h2f,8'h35,8'h1b,8'h24,8'h2c,8'h23,8'h2d,8'h2a,8'h17,8'h24,8'h27,8'h30,8'h2b,8'h26,8'h19,8'h40,8'hb6,8'hf9,8'hff,8'hc2,8'h60,8'h74,8'h7d,8'h7e,8'h79,8'h5a,8'h3f,8'hc9,8'hff,8'hff,8'hff,8'hff,8'hf7,8'hda,8'hd4,8'hd4,8'hce,8'hcc,8'hcb,8'hc6,8'hc3,8'hb9,8'h72,8'h53,8'h76,8'h72,8'h71,8'h70,8'h6e,8'h6e,8'h6a,8'h6c,8'h6e,8'h73,8'h7d,8'h7a,8'h7b,8'h79,8'h4d,8'h79,8'hfd,8'hf6,8'h72,8'h20,8'h1d,8'h2a,8'h2f,8'hbe,8'hff,8'hc0,8'h50,8'h80,8'h86,8'h85,8'h86,8'h83,8'h84,8'h85,8'h67,8'h76,8'hff,8'hff,8'hff,8'hfb,8'hf4,8'hf2,8'hee,8'he6,8'hd4,8'hc7,8'hbd,8'had,8'h81,8'h44,8'h5f,8'h81,8'h74,8'h71,8'h70,8'h6e,8'h6f,8'h75,8'h71,8'h74,8'h64,8'h2c,8'h42,8'h4f,8'h69,8'h54,8'hb2,8'hff,8'hed,8'h5d,8'h17,8'h1f,8'h22,8'h28,8'h88,8'hfa,8'hff,8'h8a,8'h3c,8'h70,8'h74,8'h6e,8'h6e,8'h71,8'h75,8'h78,8'h75,8'h72,8'h77,8'h6d,8'h62,8'h5c,8'h44,8'h4f,8'h70,8'h71,8'h72,8'h70,8'h70,8'h6f,8'h64,8'h3f,8'hb3,8'hff,8'hb3,8'h42,8'h98,8'hd1,8'hd4,8'he0,8'heb,8'hf6,8'hfb,8'hfa,8'hec,8'he5,8'hdd,8'hcd,8'hc6,8'hb5,8'h91,8'h76,8'h51,8'h4e,8'h68,8'h67,8'h6a,8'h68,8'h6c,8'h68,8'h6a,8'h69,8'h6a,8'h6c,8'h6d,8'h72,8'h77,8'h88,8'h5a,8'h5b,8'hf0,8'hff,8'h88,8'h2a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h31,8'ha1,8'hfc,8'hee,8'h6e,8'h6d,8'h82,8'h7e,8'h7b,8'h7f,8'h7a,8'h7e,8'h67,8'h5d,8'hdb,8'hff,8'hef,8'h7f,8'h3e,8'h2b,8'h24,8'h21,8'h23,8'h20,8'h14,8'h10,8'h21,8'h25,8'h22,8'h16,8'h1f,8'h20,8'h2a,8'h30,8'h47,8'h22,8'h0f,8'h4c,8'hd2,8'hff,8'hee,8'h73,8'h68,8'h79,8'h7e,8'h7e,8'h67,8'h4b,8'hd6,8'hff,8'hf9,8'hfa,8'hf4,8'hf2,8'hf1,8'hf7,8'hf4,8'hf9,8'hff,8'hff,8'hfd,8'hfb,8'hff,8'hbc,8'h3d,8'h6e,8'h71,8'h6c,8'h6d,8'h6e,8'h71,8'h74,8'h6e,8'h6e,8'h73,8'h75,8'h74,8'h75,8'h73,8'h4b,8'h8a,8'hff,8'hf2,8'h69,8'h1a,8'h20,8'h2a,8'h33,8'hc6,8'hff,8'ha5,8'h4a,8'h7e,8'h82,8'h83,8'h83,8'h81,8'h83,8'h86,8'h6c,8'h7a,8'hff,8'hfc,8'hd4,8'hc0,8'hca,8'hd4,8'hed,8'hf9,8'hff,8'hff,8'hff,8'hfe,8'hfd,8'h92,8'h39,8'h83,8'h78,8'h72,8'h74,8'h73,8'h72,8'h73,8'h79,8'h71,8'h30,8'h25,8'h60,8'h7c,8'h7a,8'h50,8'hc1,8'hff,8'he1,8'h4b,8'h3d,8'h33,8'h04,8'h29,8'hc2,8'hff,8'hef,8'h63,8'h52,8'h6f,8'h6d,8'h76,8'h79,8'h78,8'h7a,8'h7d,8'h7d,8'h75,8'h58,8'h3e,8'h45,8'h4f,8'h24,8'h53,8'h7d,8'h73,8'h6f,8'h70,8'h73,8'h77,8'h61,8'h4a,8'hc9,8'hff,8'ha2,8'h2b,8'h31,8'h3e,8'h40,8'h4c,8'h63,8'h70,8'h8d,8'haa,8'hca,8'he1,8'hea,8'hf8,8'hff,8'hfc,8'hf2,8'hef,8'hcf,8'h53,8'h5b,8'h69,8'h68,8'h69,8'h68,8'h63,8'h67,8'h6e,8'h70,8'h70,8'h6f,8'h77,8'h78,8'h7c,8'h5a,8'h58,8'hee,8'hff,8'h88,8'h2a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h5e,8'he3,8'hff,8'hb1,8'h41,8'h76,8'h78,8'h77,8'h7a,8'h79,8'h7e,8'h79,8'h56,8'h6c,8'hf3,8'hff,8'he1,8'h59,8'h37,8'h40,8'h2d,8'h1f,8'h22,8'h20,8'h07,8'h1d,8'h20,8'h13,8'h10,8'h11,8'h04,8'h12,8'h10,8'h1f,8'h26,8'h23,8'h1c,8'h28,8'ha5,8'hff,8'hf8,8'h7f,8'h62,8'h82,8'h7c,8'h7f,8'h81,8'h56,8'h94,8'hff,8'hfe,8'heb,8'h97,8'h74,8'h70,8'h75,8'h95,8'hd7,8'hf8,8'hf8,8'hfe,8'hff,8'he4,8'h79,8'h44,8'h72,8'h6d,8'h69,8'h67,8'h6c,8'h6e,8'h72,8'h73,8'h76,8'h76,8'h77,8'h75,8'h74,8'h73,8'h4d,8'h94,8'hff,8'hed,8'h65,8'h20,8'h21,8'h2a,8'h3a,8'hcc,8'hff,8'h9b,8'h53,8'h7e,8'h7d,8'h7d,8'h7d,8'h7d,8'h81,8'h89,8'h6a,8'h7c,8'hff,8'hed,8'h67,8'h33,8'h34,8'h41,8'h80,8'hc0,8'hf8,8'hfa,8'hfd,8'hff,8'hf1,8'h7a,8'h3e,8'h80,8'h79,8'h76,8'h77,8'h7a,8'h78,8'h7e,8'h7c,8'h62,8'h34,8'h67,8'h7d,8'h7c,8'h71,8'h4a,8'hc2,8'hff,8'hd5,8'h3b,8'h27,8'h1f,8'h00,8'h48,8'hdf,8'hff,8'hd5,8'h53,8'h66,8'h74,8'h73,8'h77,8'h7a,8'h7c,8'h7f,8'h75,8'h58,8'h3f,8'h49,8'h82,8'hcb,8'hb1,8'h38,8'h61,8'h7b,8'h72,8'h70,8'h73,8'h75,8'h6e,8'h4d,8'h51,8'he3,8'hfb,8'h8a,8'h24,8'h34,8'h25,8'h14,8'h19,8'h0b,8'h0f,8'h28,8'h2b,8'h34,8'h49,8'h6e,8'hdb,8'hfc,8'hfa,8'hfb,8'hff,8'he1,8'h4a,8'h59,8'h68,8'h67,8'h66,8'h69,8'h65,8'h64,8'h6f,8'h70,8'h71,8'h74,8'h78,8'h78,8'h80,8'h58,8'h5e,8'hf1,8'hff,8'h89,8'h2a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h38,8'hb1,8'hff,8'hf5,8'h60,8'h4f,8'h7a,8'h74,8'h7b,8'h79,8'h78,8'h82,8'h7a,8'h55,8'h82,8'hff,8'hff,8'hc9,8'h42,8'h17,8'h3d,8'h3f,8'h44,8'h24,8'h17,8'h14,8'h21,8'h1f,8'h1d,8'h17,8'h11,8'h07,8'h16,8'h16,8'h14,8'h1c,8'h24,8'h23,8'h24,8'h96,8'hfc,8'hf7,8'h80,8'h5f,8'h82,8'h7a,8'h7e,8'h83,8'h65,8'h64,8'hec,8'hff,8'hec,8'h7b,8'h32,8'h1f,8'h38,8'hb6,8'hec,8'hfc,8'hff,8'hea,8'ha4,8'h5f,8'h3a,8'h67,8'h76,8'h6d,8'h70,8'h71,8'h6e,8'h6d,8'h72,8'h73,8'h75,8'h79,8'h76,8'h75,8'h75,8'h79,8'h4e,8'h94,8'hff,8'hea,8'h65,8'h23,8'h25,8'h22,8'h35,8'hce,8'hff,8'h97,8'h52,8'h7d,8'h7d,8'h7a,8'h81,8'h7f,8'h81,8'h88,8'h6e,8'h7d,8'hff,8'hea,8'h52,8'h25,8'h26,8'h26,8'h28,8'h78,8'hf7,8'hff,8'hf4,8'hc2,8'h6b,8'h39,8'h61,8'h81,8'h7a,8'h79,8'h77,8'h77,8'h7d,8'h7f,8'h7e,8'h79,8'h75,8'h83,8'h7f,8'h80,8'h6f,8'h46,8'hc3,8'hff,8'hcd,8'h35,8'h04,8'h0f,8'h07,8'h66,8'hef,8'hff,8'hb2,8'h48,8'h71,8'h7b,8'h7e,8'h77,8'h7a,8'h74,8'h57,8'h48,8'h5e,8'h94,8'hd9,8'hfa,8'hff,8'ha3,8'h35,8'h6a,8'h74,8'h72,8'h6e,8'h71,8'h70,8'h6e,8'h44,8'h68,8'hf3,8'hf0,8'h6d,8'h18,8'h2b,8'h22,8'h12,8'h19,8'h14,8'h08,8'h29,8'h39,8'h1d,8'h21,8'h72,8'heb,8'hfe,8'hff,8'hfc,8'hd0,8'h6b,8'h35,8'h69,8'h68,8'h65,8'h66,8'h67,8'h6c,8'h65,8'h66,8'h72,8'h6e,8'h71,8'h7a,8'h7a,8'h86,8'h57,8'h66,8'hf6,8'hff,8'h8a,8'h2a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h5b,8'he7,8'hff,8'hc6,8'h38,8'h6c,8'h75,8'h73,8'h77,8'h7a,8'h77,8'h7b,8'h76,8'h52,8'ha6,8'hff,8'hfc,8'hb2,8'h32,8'h23,8'h2b,8'h2d,8'h44,8'h23,8'h18,8'h30,8'h46,8'h20,8'h1f,8'h18,8'h1c,8'h14,8'h17,8'h1e,8'h1f,8'h2a,8'h40,8'h3b,8'h37,8'haf,8'hfe,8'hf0,8'h71,8'h60,8'h7f,8'h7e,8'h80,8'h80,8'h76,8'h53,8'hb6,8'hff,8'hf8,8'hba,8'h52,8'h0e,8'h5e,8'hf1,8'hff,8'hff,8'hc2,8'h63,8'h42,8'h52,8'h68,8'h72,8'h6c,8'h6e,8'h77,8'h77,8'h70,8'h70,8'h60,8'h68,8'h7d,8'h7a,8'h7a,8'h7e,8'h7e,8'h82,8'h4f,8'h96,8'hff,8'heb,8'h7b,8'h38,8'h2e,8'h33,8'h40,8'hd2,8'hff,8'h94,8'h58,8'h82,8'h81,8'h83,8'h83,8'h84,8'h86,8'h8f,8'h6f,8'h7d,8'hff,8'hea,8'h52,8'h25,8'h26,8'h26,8'h3c,8'hb8,8'hf9,8'hc6,8'h67,8'h38,8'h3d,8'h65,8'h7b,8'h7f,8'h81,8'h7f,8'h75,8'h67,8'h52,8'h42,8'h74,8'h8b,8'h83,8'h84,8'h88,8'h87,8'h74,8'h51,8'hca,8'hff,8'hc8,8'h36,8'h0c,8'h1a,8'h0d,8'h71,8'hf5,8'hff,8'h8a,8'h4e,8'h7d,8'h81,8'h85,8'h85,8'h77,8'h48,8'h50,8'h98,8'he3,8'hfc,8'hfe,8'hfa,8'hfd,8'h88,8'h3f,8'h74,8'h77,8'h7d,8'h77,8'h76,8'h77,8'h6b,8'h34,8'h80,8'hfe,8'he4,8'h52,8'h15,8'h15,8'h12,8'h1b,8'h14,8'h1c,8'h1f,8'h26,8'h44,8'h27,8'h52,8'hd8,8'hfd,8'hff,8'he6,8'h86,8'h3c,8'h35,8'h63,8'h71,8'h70,8'h70,8'h6f,8'h72,8'h61,8'h3f,8'h39,8'h6d,8'h75,8'h77,8'h78,8'h76,8'h81,8'h5c,8'h6f,8'hf9,8'hff,8'h8a,8'h2a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h2c,8'h9a,8'hfc,8'hfb,8'h77,8'h40,8'h7c,8'h75,8'h7d,8'h75,8'h75,8'h73,8'h7a,8'h72,8'h52,8'hc1,8'hff,8'hfa,8'h9f,8'h32,8'h33,8'h24,8'h2a,8'h36,8'h21,8'h1c,8'h23,8'h24,8'h1f,8'h22,8'h1c,8'h1f,8'h1d,8'h1d,8'h1e,8'h20,8'h31,8'h32,8'h38,8'h6f,8'he2,8'hff,8'hdd,8'h5b,8'h67,8'h7e,8'h80,8'h82,8'h83,8'h85,8'h5f,8'h81,8'hf9,8'hff,8'hd8,8'h5d,8'h13,8'h6d,8'hf5,8'hff,8'hcc,8'h57,8'h54,8'h74,8'h81,8'h81,8'h7a,8'h7e,8'h7b,8'h7c,8'h79,8'h60,8'h48,8'h2a,8'h55,8'h89,8'h7f,8'h7e,8'h86,8'h86,8'h81,8'h43,8'h92,8'hff,8'heb,8'h72,8'h38,8'h30,8'h38,8'h42,8'hda,8'hff,8'h91,8'h50,8'h7e,8'h7f,8'h85,8'h84,8'h85,8'h84,8'h8a,8'h71,8'h7c,8'hff,8'he8,8'h52,8'h25,8'h26,8'h27,8'h71,8'hee,8'hba,8'h38,8'h2e,8'h63,8'h7e,8'h84,8'h80,8'h79,8'h75,8'h75,8'h5d,8'h39,8'h31,8'h22,8'h5d,8'h75,8'h6d,8'h72,8'h73,8'h6f,8'h57,8'h5e,8'he2,8'hff,8'hcc,8'h42,8'h1f,8'h14,8'h0d,8'h82,8'hfb,8'hf9,8'h67,8'h3d,8'h5f,8'h61,8'h61,8'h63,8'h48,8'h3d,8'hbe,8'hf9,8'hfb,8'he9,8'he5,8'hf6,8'hfc,8'h73,8'h30,8'h50,8'h53,8'h5a,8'h55,8'h4e,8'h52,8'h41,8'h2e,8'hac,8'hff,8'hcb,8'h37,8'h0f,8'h0f,8'h13,8'h19,8'h0c,8'h17,8'h1d,8'h1e,8'h37,8'h27,8'h98,8'hfb,8'hff,8'hc6,8'h4e,8'h16,8'h18,8'h2e,8'h37,8'h31,8'h32,8'h30,8'h2f,8'h2f,8'h34,8'h35,8'h23,8'h2d,8'h2c,8'h30,8'h2f,8'h2f,8'h33,8'h27,8'h6f,8'hfa,8'hff,8'h8a,8'h2a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h25,8'h49,8'hd8,8'hff,8'hdb,8'h3f,8'h4a,8'h64,8'h63,8'h67,8'h6a,8'h67,8'h68,8'h68,8'h5c,8'h4f,8'hdc,8'hff,8'hf5,8'h96,8'h31,8'h31,8'h25,8'h22,8'h20,8'h1f,8'h20,8'h1a,8'h1b,8'h22,8'h22,8'h20,8'h20,8'h1f,8'h21,8'h2d,8'h23,8'h17,8'h20,8'h53,8'hc5,8'hfc,8'hf9,8'h95,8'h37,8'h54,8'h55,8'h54,8'h55,8'h54,8'h52,8'h42,8'h42,8'hcc,8'hff,8'hf4,8'ha4,8'h30,8'h7c,8'hfa,8'hfe,8'h77,8'h30,8'h4f,8'h4e,8'h52,8'h51,8'h4b,8'h49,8'h4a,8'h4b,8'h50,8'h61,8'h6d,8'h49,8'h2c,8'h40,8'h46,8'h4b,8'h4a,8'h42,8'h3d,8'h29,8'h97,8'hff,8'heb,8'h62,8'h0e,8'h1d,8'h0d,8'h45,8'he2,8'hff,8'h8f,8'h29,8'h2e,8'h2a,8'h28,8'h2d,8'h2d,8'h2a,8'h2d,8'h27,8'h76,8'hff,8'he8,8'h52,8'h25,8'h26,8'h2a,8'ha9,8'he9,8'h55,8'h02,8'h21,8'h2b,8'h2d,8'h25,8'h20,8'h26,8'h28,8'h3b,8'h58,8'h96,8'hae,8'h36,8'h0d,8'h14,8'h0e,8'h01,8'h07,8'h1a,8'h09,8'h4a,8'hec,8'hff,8'hc9,8'h61,8'h29,8'h0d,8'h1e,8'ha0,8'hff,8'he7,8'h3d,8'h00,8'h00,8'h00,8'h04,8'h01,8'h0a,8'h68,8'hf9,8'hf4,8'hbd,8'h7f,8'h99,8'he8,8'hde,8'h47,8'h07,8'h04,8'h00,8'h00,8'h00,8'h00,8'h12,8'h0c,8'h46,8'he4,8'hfe,8'h9c,8'h27,8'h11,8'h14,8'h14,8'h29,8'h27,8'h12,8'h05,8'h18,8'h2b,8'h46,8'hd5,8'hff,8'hd9,8'h44,8'h0c,8'h03,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0b,8'h31,8'h57,8'h9d,8'h98,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'h15,8'h7a,8'hff,8'hff,8'h8b,8'h2a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h78,8'hef,8'hff,8'h90,8'h20,8'h18,8'h17,8'h14,8'h17,8'h11,8'h0d,8'h17,8'h21,8'h0b,8'h42,8'he6,8'hff,8'hef,8'h9a,8'h31,8'h1f,8'h20,8'h1a,8'h10,8'h1f,8'h20,8'h20,8'h1f,8'h10,8'h16,8'h1b,8'h22,8'h28,8'h39,8'h4b,8'h40,8'h32,8'h79,8'hdc,8'hf7,8'hf8,8'ha8,8'h2a,8'h02,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h7c,8'hff,8'hff,8'hd2,8'h52,8'ha3,8'hff,8'hf0,8'h58,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h18,8'h51,8'h98,8'he1,8'hf0,8'h71,8'h0e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h16,8'ha1,8'hff,8'he8,8'h6a,8'h27,8'h22,8'h1f,8'h50,8'he9,8'hff,8'h8a,8'h07,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h73,8'hff,8'hea,8'h52,8'h25,8'h25,8'h37,8'hc6,8'hcc,8'h2d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h4b,8'hb5,8'hed,8'hff,8'hd8,8'h39,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h4c,8'hee,8'hff,8'hb3,8'h4c,8'h32,8'h10,8'h2d,8'hc3,8'hff,8'hc7,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0e,8'h94,8'hff,8'hef,8'hb1,8'hb8,8'he4,8'hc5,8'h55,8'h0a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1d,8'h95,8'hff,8'he9,8'h61,8'h20,8'h20,8'h1f,8'h13,8'h1e,8'h20,8'h20,8'h15,8'h1f,8'h30,8'h6f,8'hf2,8'hff,8'h97,8'h16,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1b,8'h5b,8'hc2,8'hf0,8'hff,8'had,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0c,8'h7f,8'hff,8'hff,8'h8b,8'h2a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h25,8'h00,8'h00},
'{8'h00,8'h00,8'h25,8'h38,8'hb8,8'hff,8'hee,8'h54,8'h1e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h43,8'he2,8'hff,8'hed,8'h79,8'h21,8'h20,8'h1f,8'h17,8'h17,8'h20,8'h21,8'h20,8'h1f,8'h28,8'h2a,8'h1a,8'h23,8'h2a,8'h38,8'h2b,8'h51,8'h96,8'he6,8'hf8,8'hf4,8'ha9,8'h2f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3c,8'hdb,8'hff,8'hf4,8'h9d,8'hc4,8'hff,8'hdf,8'h3f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h4b,8'hd4,8'hff,8'hff,8'hf0,8'h56,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1d,8'haf,8'hff,8'he8,8'h62,8'h1e,8'h1f,8'h20,8'h5a,8'hec,8'hff,8'h8a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h75,8'hff,8'heb,8'h53,8'h25,8'h25,8'h4c,8'hdf,8'hbc,8'h1f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2f,8'hc0,8'hff,8'hff,8'hff,8'hd3,8'h34,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h4b,8'hf0,8'hff,8'ha9,8'h2b,8'h34,8'h13,8'h5a,8'he6,8'hff,8'ha0,8'h0c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h18,8'hb0,8'hff,8'hfd,8'hed,8'hca,8'h7f,8'h33,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3c,8'hdd,8'hff,8'hc8,8'h50,8'h1f,8'h10,8'h0c,8'h14,8'h1f,8'h18,8'h23,8'h32,8'h15,8'h1e,8'h84,8'hfd,8'hfe,8'h7c,8'h13,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h5f,8'he0,8'hff,8'hfd,8'hff,8'ha0,8'h12,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h08,8'h80,8'hff,8'hff,8'h8b,8'h2a,8'h00,8'h00,8'h00,8'h00,8'h27,8'h2a,8'h3c,8'h61,8'h7f,8'h5a,8'h2a,8'h00},
'{8'h00,8'h00,8'h25,8'h62,8'he4,8'hff,8'hc0,8'h2c,8'h0e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h37,8'hd3,8'hff,8'hf6,8'h91,8'h23,8'h1f,8'h22,8'h20,8'h1f,8'h20,8'h20,8'h1f,8'h23,8'h33,8'h2f,8'h25,8'h2e,8'h23,8'h3a,8'h74,8'hbe,8'hef,8'hff,8'hd4,8'h83,8'h31,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h11,8'h89,8'hff,8'hff,8'he4,8'hea,8'hff,8'hc2,8'h2a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2a,8'haa,8'hff,8'hf2,8'hf2,8'he9,8'h46,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'hbe,8'hff,8'hea,8'h62,8'h1d,8'h3a,8'h66,8'hae,8'hf9,8'hff,8'h86,8'h06,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h77,8'hff,8'heb,8'h52,8'h25,8'h25,8'h63,8'he8,8'h8f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h64,8'hf7,8'hf6,8'hb6,8'he3,8'hc9,8'h31,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h61,8'hf8,8'hff,8'h96,8'h20,8'h25,8'h3f,8'haf,8'hfd,8'hff,8'h7d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0f,8'h69,8'h8b,8'h81,8'h50,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h28,8'h6b,8'hbe,8'hff,8'hea,8'h77,8'h44,8'h27,8'h1a,8'h0b,8'h13,8'h17,8'h14,8'h1d,8'h1c,8'h16,8'h21,8'ha4,8'hff,8'hf0,8'h5c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'had,8'hff,8'hd8,8'hca,8'hfc,8'h97,8'h08,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h06,8'h7f,8'hff,8'hff,8'h88,8'h28,8'h00,8'h2e,8'h42,8'h64,8'h81,8'h95,8'hca,8'hea,8'hee,8'h88,8'h2a,8'h25},
'{8'h00,8'h25,8'h28,8'h88,8'hf8,8'hff,8'h80,8'h12,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'ha5,8'hff,8'hff,8'hcd,8'h51,8'h20,8'h1f,8'h21,8'h20,8'h1e,8'h1e,8'h1f,8'h22,8'h21,8'h1d,8'h27,8'h43,8'h61,8'hb1,8'hee,8'hff,8'hfb,8'hc0,8'h4d,8'h02,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h41,8'he1,8'hff,8'hfa,8'hfc,8'hff,8'ha6,8'h17,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h43,8'hdd,8'hfd,8'ha6,8'hb7,8'he0,8'h3c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2d,8'hc8,8'hff,8'he3,8'h75,8'h7f,8'hc9,8'hf0,8'hfb,8'hff,8'hff,8'h80,8'h08,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h75,8'hff,8'hea,8'h53,8'h26,8'h24,8'h7e,8'hee,8'h6c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h95,8'hff,8'hd1,8'h58,8'hc8,8'hbd,8'h2a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h79,8'hff,8'hff,8'h9c,8'h48,8'h7a,8'hcc,8'hf5,8'hfe,8'hf6,8'h4e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h08,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h58,8'hb8,8'hf9,8'hff,8'hf2,8'h96,8'h2c,8'h1b,8'h3c,8'h2b,8'h11,8'h12,8'h0c,8'h28,8'h38,8'h26,8'h2c,8'h2d,8'hbc,8'hff,8'he1,8'h3e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3c,8'hcf,8'hff,8'h8e,8'h86,8'hf3,8'h8b,8'h11,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0b,8'h80,8'hff,8'hff,8'h9e,8'h4a,8'h6f,8'h9c,8'hd4,8'hf2,8'hff,8'hff,8'hff,8'hff,8'hbc,8'h44,8'h25,8'h00},
'{8'h00,8'h25,8'h40,8'hc0,8'hff,8'hef,8'h4e,8'h0f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h14,8'h6c,8'hf4,8'hff,8'hf6,8'hc5,8'h6b,8'h3b,8'h31,8'h2b,8'h27,8'h2a,8'h2c,8'h31,8'h34,8'h43,8'h66,8'ha1,8'hdf,8'hf7,8'hfe,8'hec,8'ha3,8'h42,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h22,8'ha3,8'hff,8'hfc,8'hfa,8'hff,8'h92,8'h0b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h5e,8'hf1,8'hf1,8'h71,8'hac,8'hc8,8'h29,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h28,8'hd6,8'hff,8'hf8,8'he7,8'hf1,8'hfc,8'hff,8'hff,8'hff,8'hff,8'h6e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h74,8'hff,8'heb,8'h53,8'h25,8'h27,8'h8c,8'he7,8'h4d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h13,8'hba,8'hff,8'he8,8'hb5,8'hec,8'h9c,8'h12,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h84,8'hff,8'hff,8'hd9,8'hcf,8'hf2,8'hfc,8'hfe,8'hff,8'hec,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h28,8'h4a,8'ha1,8'heb,8'hff,8'hfa,8'hdd,8'h8f,8'h38,8'h1d,8'h16,8'h12,8'h17,8'h1c,8'h13,8'h0e,8'h26,8'h2a,8'h35,8'h4f,8'h4f,8'hd5,8'hff,8'hd0,8'h2f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h4e,8'he7,8'hfd,8'hc3,8'hd8,8'hf5,8'h69,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0e,8'h85,8'hff,8'hff,8'he5,8'hd0,8'hf6,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfd,8'hc6,8'h50,8'h00,8'h00,8'h00},
'{8'h00,8'h27,8'h6c,8'hea,8'hff,8'hcd,8'h2e,8'h18,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2f,8'h9a,8'hfe,8'hff,8'hfb,8'he4,8'hc5,8'hba,8'hac,8'ha5,8'ha4,8'ha6,8'hb3,8'hbc,8'hcf,8'he6,8'hf8,8'hff,8'he7,8'ha7,8'h5a,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h53,8'hec,8'hff,8'hfc,8'hf9,8'h6e,8'h03,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6e,8'hf8,8'hf5,8'hc7,8'hec,8'hb5,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2a,8'hdc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hf8,8'hcc,8'he5,8'hfa,8'h62,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h76,8'hff,8'heb,8'h53,8'h25,8'h32,8'haf,8'hd4,8'h30,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2c,8'hd7,8'hff,8'hfc,8'hff,8'hde,8'h4c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8c,8'hff,8'hff,8'hfb,8'hfc,8'hff,8'hff,8'he4,8'he8,8'hca,8'h29,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1f,8'h72,8'hbf,8'he0,8'hff,8'hfe,8'hdc,8'h92,8'h56,8'h2c,8'h20,8'h22,8'h1b,8'h0e,8'h16,8'h18,8'h10,8'h1e,8'h2c,8'h2e,8'h2f,8'h26,8'h5f,8'he5,8'hff,8'hb0,8'h21,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h5b,8'hf0,8'hff,8'hff,8'hfb,8'hb5,8'h31,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h06,8'h84,8'hff,8'hff,8'hff,8'hff,8'hf2,8'hbd,8'hb5,8'hf6,8'hff,8'hfd,8'hbd,8'h4c,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h2c,8'h92,8'hf9,8'hff,8'h9a,8'h21,8'h0b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2a,8'h8e,8'hed,8'hff,8'hff,8'hfd,8'hfc,8'hfa,8'hf8,8'hf9,8'hfb,8'hfe,8'hfe,8'hff,8'hff,8'hec,8'ha6,8'h4c,8'h15,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'hab,8'hff,8'hff,8'hf0,8'h52,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8a,8'hfb,8'hf9,8'hff,8'hf8,8'h79,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h30,8'hde,8'hff,8'hff,8'hff,8'hf8,8'hc0,8'h68,8'h68,8'he1,8'hf6,8'h5a,8'h02,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h76,8'hff,8'hec,8'h53,8'h24,8'h39,8'hc1,8'haf,8'h23,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h42,8'hea,8'hff,8'hfc,8'hdc,8'h64,8'h02,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8c,8'hff,8'hff,8'hff,8'hfe,8'he1,8'h8a,8'h49,8'ha4,8'hb3,8'h21,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0b,8'h71,8'hef,8'hff,8'hfe,8'he6,8'ha1,8'h52,8'h44,8'h39,8'h20,8'h20,8'h1f,8'h1e,8'h1f,8'h1b,8'h18,8'h13,8'h20,8'h38,8'h43,8'h3f,8'h2a,8'h6b,8'hf1,8'hff,8'h8d,8'h11,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h84,8'hfe,8'hff,8'hf0,8'h96,8'h33,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h02,8'h87,8'hff,8'hff,8'he9,8'ha8,8'h54,8'h30,8'h94,8'hfe,8'hff,8'hc1,8'h4a,8'h25,8'h00,8'h00,8'h00,8'h00},
'{8'h25,8'h32,8'hb8,8'hff,8'hff,8'h77,8'h0c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h22,8'h63,8'hc1,8'he4,8'hf1,8'hf8,8'hf7,8'hf5,8'hf5,8'hf0,8'he8,8'hdc,8'hcf,8'ha2,8'h59,8'h1a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h5f,8'hef,8'hff,8'he8,8'h49,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h92,8'hec,8'hdc,8'hd5,8'h92,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h28,8'ha9,8'hdf,8'hd9,8'hab,8'h64,8'h33,8'h59,8'hcf,8'hff,8'hf3,8'h54,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h75,8'hff,8'hed,8'h53,8'h24,8'h4e,8'hd9,8'h90,8'h15,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h31,8'hbc,8'hc8,8'h85,8'h3b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h62,8'he5,8'hea,8'hcd,8'h87,8'h3e,8'h2a,8'h6a,8'he2,8'ha3,8'h21,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'h00,8'h00,8'h00,8'h43,8'hd6,8'hff,8'hea,8'hb1,8'h63,8'h34,8'h2b,8'h4c,8'h56,8'h42,8'h43,8'h1f,8'h16,8'h20,8'h2a,8'h1f,8'h0f,8'h15,8'h20,8'h34,8'h2a,8'h31,8'h86,8'hfb,8'hf8,8'h68,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h80,8'hdd,8'hba,8'h5d,8'h1a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h06,8'h6e,8'hc9,8'h92,8'h46,8'h1f,8'h27,8'h83,8'hf0,8'hff,8'hca,8'h54,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h25,8'h37,8'hcc,8'hff,8'hf6,8'h5a,8'h0a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2d,8'h47,8'h65,8'h71,8'h72,8'h70,8'h6d,8'h66,8'h53,8'h3d,8'h2c,8'h05,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'hae,8'hff,8'hd0,8'h2c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h39,8'h59,8'h3c,8'h2a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h29,8'h36,8'h33,8'h23,8'h24,8'h77,8'he5,8'hff,8'hff,8'hee,8'h4e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h76,8'hff,8'hed,8'h54,8'h23,8'h5d,8'hdd,8'h69,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2e,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h53,8'h4b,8'h2f,8'h0a,8'h29,8'h9e,8'hf1,8'hff,8'h80,8'h10,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h29,8'h56,8'h88,8'h4e,8'h01,8'h00,8'h1f,8'h9d,8'hff,8'hfc,8'hc5,8'h7b,8'h6c,8'h7f,8'h8d,8'h95,8'h98,8'h9d,8'h92,8'h7a,8'h5c,8'h55,8'h77,8'h34,8'h1e,8'h28,8'h1c,8'h22,8'h1f,8'h26,8'hac,8'hff,8'hec,8'h4d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h28,8'h41,8'h29,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h21,8'h2d,8'h1d,8'h14,8'h2d,8'ha1,8'hf7,8'hff,8'hbf,8'h4e,8'h28,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h25,8'h3c,8'he3,8'hff,8'he9,8'h40,8'h08,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h72,8'hfd,8'haf,8'h1d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h85,8'hf2,8'hff,8'hff,8'hff,8'hed,8'h4a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h76,8'hff,8'hec,8'h53,8'h26,8'h7c,8'he1,8'h4a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2e,8'h9e,8'hfc,8'hff,8'hfe,8'h6d,8'h07,8'h00,8'h00,8'h00,8'h01,8'h21,8'h39,8'h6c,8'hb8,8'heb,8'he9,8'h58,8'h04,8'h00,8'h47,8'he3,8'hff,8'hfb,8'hec,8'he5,8'he9,8'hf1,8'hf6,8'hf8,8'hf7,8'hf6,8'hf2,8'hee,8'he0,8'hcf,8'hc2,8'h80,8'h71,8'h52,8'h26,8'h1c,8'h19,8'h36,8'hc6,8'hff,8'hda,8'h33,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h08,8'h25,8'h8c,8'hfa,8'hff,8'hc8,8'h4d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h25,8'h3f,8'heb,8'hff,8'he6,8'h34,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h05,8'h2f,8'h5a,8'haa,8'hfc,8'h89,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h36,8'h98,8'hf7,8'hff,8'he3,8'hc2,8'hf7,8'hed,8'h48,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h73,8'hff,8'hee,8'h52,8'h31,8'hac,8'hd0,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'h46,8'hac,8'hff,8'hff,8'hff,8'hff,8'h79,8'h23,8'h26,8'h3c,8'h60,8'h6c,8'ha0,8'hd7,8'hf3,8'hff,8'hfb,8'h93,8'h23,8'h00,8'h01,8'h81,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hff,8'hff,8'hfd,8'hf6,8'hea,8'hd3,8'h9a,8'h59,8'h25,8'h16,8'h4a,8'hde,8'hff,8'hc2,8'h2a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h14,8'h32,8'h8c,8'hf2,8'hff,8'hc9,8'h56,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h25,8'h3f,8'hec,8'hff,8'he4,8'h30,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2c,8'h67,8'hb9,8'hf3,8'hff,8'hfd,8'h6a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3e,8'hbb,8'hff,8'hff,8'hd3,8'h65,8'h42,8'hd7,8'hee,8'h49,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h09,8'h85,8'hff,8'hec,8'h50,8'h51,8'he8,8'hb0,8'h28,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h4f,8'hd2,8'hff,8'hfd,8'hea,8'hff,8'hff,8'hd7,8'ha4,8'hbd,8'he1,8'hf8,8'hf9,8'hfc,8'hfe,8'hfe,8'hff,8'haf,8'h2b,8'h00,8'h00,8'h25,8'ha7,8'hff,8'hff,8'hf0,8'hd7,8'hc9,8'hb9,8'ha4,8'ha0,8'ha0,8'ha7,8'hbc,8'hd0,8'he6,8'hfc,8'hff,8'hff,8'hff,8'hfe,8'hf7,8'hd8,8'h77,8'h28,8'h62,8'hec,8'hff,8'h97,8'h0d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0f,8'h2e,8'haa,8'hfe,8'hff,8'hc9,8'h4f,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h25,8'h3d,8'he6,8'hff,8'he6,8'h37,8'h0a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h61,8'hb1,8'hf1,8'hff,8'hff,8'hff,8'hed,8'h48,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h45,8'hb7,8'hff,8'hff,8'hcf,8'h58,8'h28,8'h33,8'hc4,8'hed,8'h4b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2d,8'hbe,8'hff,8'he3,8'h4b,8'h68,8'hf0,8'h89,8'h0b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h18,8'h5c,8'hd5,8'hff,8'hfa,8'had,8'h7d,8'hea,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hfb,8'hf6,8'hf2,8'hf8,8'hfe,8'hea,8'h56,8'h0b,8'h00,8'h00,8'h0b,8'h5b,8'h9a,8'h8d,8'h63,8'h39,8'h28,8'h22,8'h1d,8'h17,8'h13,8'h11,8'h22,8'h2f,8'h46,8'h72,8'hb5,8'hec,8'hff,8'hff,8'hff,8'hfa,8'he5,8'h88,8'h98,8'hf8,8'hff,8'h7d,8'h0c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h09,8'h2f,8'h30,8'h06,8'h00,8'h00,8'h00,8'h00,8'h00,8'h28,8'h92,8'hf9,8'hff,8'hcb,8'h57,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h25,8'h37,8'hce,8'hff,8'hf3,8'h57,8'h1d,8'h05,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h30,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h06,8'h3b,8'h81,8'hb6,8'hec,8'hff,8'hff,8'hf2,8'hd9,8'hf2,8'he6,8'h34,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h4a,8'h7d,8'h2d,8'h00,8'h00,8'h00,8'h00,8'h09,8'h5f,8'hcd,8'hff,8'hff,8'hb5,8'h52,8'h28,8'h27,8'h40,8'hde,8'hea,8'h48,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h28,8'h94,8'hf6,8'hff,8'hb4,8'h3b,8'h8b,8'hf8,8'h75,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0e,8'h4d,8'h80,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'h22,8'h76,8'he2,8'hff,8'he2,8'h91,8'h41,8'h34,8'h88,8'hc2,8'hdc,8'hd6,8'hbe,8'h9a,8'h88,8'h83,8'h9d,8'hea,8'hfa,8'h8a,8'h1f,8'h04,8'h00,8'h06,8'h19,8'h1f,8'h1f,8'h1f,8'h13,8'h07,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h23,8'h4f,8'h81,8'hcc,8'hff,8'hff,8'hff,8'hec,8'he7,8'hfc,8'hf6,8'h58,8'h09,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h2e,8'h79,8'hc1,8'h93,8'h22,8'h00,8'h00,8'h00,8'h0b,8'h34,8'ha1,8'hf3,8'hfb,8'hbd,8'h53,8'h28,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h25,8'h31,8'hb0,8'hfe,8'hff,8'h7e,8'h11,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h28,8'h7c,8'had,8'h38,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h09,8'h33,8'h76,8'hd2,8'hfe,8'hff,8'hff,8'hf6,8'hc1,8'h68,8'h5d,8'hd5,8'he1,8'h31,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h29,8'h69,8'hda,8'he4,8'h45,8'h00,8'h00,8'h00,8'h1d,8'h6b,8'he3,8'hff,8'hf9,8'hc2,8'h49,8'h26,8'h27,8'h27,8'h43,8'he5,8'he6,8'h44,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h23,8'h8e,8'hf7,8'hff,8'hec,8'h68,8'h2a,8'h96,8'hfa,8'h71,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h16,8'h39,8'h90,8'he5,8'heb,8'h50,8'h00,8'h00,8'h00,8'h00,8'h29,8'h82,8'hf2,8'hff,8'he3,8'h70,8'h2d,8'h26,8'h00,8'h2d,8'h3a,8'h48,8'h45,8'h39,8'h2e,8'h29,8'h2f,8'h91,8'hfc,8'hd0,8'h2c,8'h12,8'h29,8'h3e,8'h56,8'h6d,8'h73,8'h73,8'h65,8'h40,8'h22,8'h0e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h05,8'h31,8'ha0,8'hf7,8'hff,8'hfd,8'hfb,8'hff,8'hf7,8'h53,8'h0e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h06,8'h29,8'h64,8'hc5,8'hfb,8'hff,8'hb6,8'h27,8'h01,8'h00,8'h16,8'h31,8'ha9,8'hff,8'hff,8'hc2,8'h4a,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h2a,8'h87,8'hf8,8'hff,8'hb7,8'h1d,8'h0a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h2a,8'h52,8'haa,8'hf7,8'hb8,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h15,8'h39,8'h73,8'hcc,8'hf9,8'hff,8'hf9,8'he0,8'hc5,8'h83,8'h40,8'h25,8'h43,8'hd0,8'he6,8'h3b,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2b,8'h44,8'h9a,8'hef,8'hff,8'hf0,8'h53,8'h07,8'h00,8'h20,8'h71,8'he4,8'hff,8'he0,8'h85,8'h3e,8'h28,8'h27,8'h27,8'h27,8'h43,8'he4,8'he3,8'h46,8'h00,8'h00,8'h00,8'h00,8'h11,8'h35,8'h92,8'hf3,8'hff,8'hef,8'h95,8'h34,8'h29,8'h94,8'hfc,8'h7c,8'h0b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h44,8'h7d,8'hd0,8'hff,8'hff,8'hfd,8'h70,8'h08,8'h00,8'h00,8'h31,8'h8c,8'hf3,8'hf5,8'hbb,8'h65,8'h2c,8'h26,8'h00,8'h00,8'h25,8'h25,8'h25,8'h25,8'h25,8'h25,8'h26,8'h5a,8'hde,8'hfa,8'h80,8'h37,8'h6b,8'had,8'he2,8'hf4,8'hfd,8'hff,8'hff,8'hfc,8'he3,8'hb3,8'h6d,8'h30,8'h21,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h87,8'hf0,8'hff,8'hfe,8'hff,8'hff,8'h86,8'h14,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h08,8'h24,8'h2d,8'h54,8'haf,8'hf2,8'hff,8'hff,8'hff,8'hbd,8'h26,8'h0b,8'h15,8'h2b,8'h91,8'hf8,8'hff,8'hc5,8'h50,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h25,8'h54,8'hd9,8'hff,8'hed,8'h52,8'h0b,8'h07,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h22,8'h50,8'ha8,8'he7,8'hff,8'hff,8'h7a,8'h0e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1d,8'h4a,8'h95,8'hcf,8'hf5,8'hff,8'hff,8'hdc,8'h85,8'h4b,8'h39,8'h29,8'h00,8'h25,8'h47,8'hd6,8'hfe,8'h7f,8'h0f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1e,8'h37,8'h6c,8'hb3,8'hda,8'hfe,8'hf5,8'hf0,8'hfb,8'h78,8'h12,8'h31,8'h94,8'heb,8'hff,8'he2,8'h60,8'h2b,8'h26,8'h27,8'h27,8'h27,8'h27,8'h43,8'he4,8'he4,8'h45,8'h00,8'h00,8'h03,8'h25,8'h6e,8'hc7,8'hfa,8'hff,8'he5,8'h77,8'h32,8'h25,8'h29,8'h7d,8'hf9,8'hbc,8'h2f,8'h00,8'h00,8'h00,8'h00,8'h04,8'h27,8'h49,8'h82,8'hbb,8'hd8,8'hf7,8'hff,8'he5,8'hdf,8'hff,8'h8c,8'h0e,8'h00,8'h42,8'hb1,8'hf4,8'hf8,8'h95,8'h38,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3c,8'hb8,8'hfe,8'hf4,8'hc3,8'hcf,8'hef,8'hfa,8'hf5,8'hf4,8'hfb,8'hfd,8'hfc,8'hff,8'hff,8'hff,8'hf4,8'hca,8'h7b,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h21,8'h7b,8'hf4,8'hff,8'hff,8'hff,8'hd5,8'h40,8'h0f,8'h0e,8'h00,8'h00,8'h0b,8'h27,8'h60,8'h95,8'hc7,8'he7,8'hff,8'hf9,8'he4,8'hef,8'hff,8'hda,8'h3e,8'h12,8'h3d,8'ha7,8'hf3,8'hfc,8'hbd,8'h4d,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h25,8'h2e,8'h9a,8'hfd,8'hff,8'hb5,8'h29,8'h11,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1a,8'h34,8'h85,8'he0,8'hff,8'hff,8'hff,8'hef,8'h56,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0d,8'h3b,8'h90,8'hdc,8'hff,8'hff,8'hff,8'he3,8'ha0,8'h59,8'h2a,8'h25,8'h25,8'h00,8'h00,8'h25,8'h3c,8'hc3,8'hff,8'he6,8'h6c,8'h24,8'h12,8'h17,8'h22,8'h32,8'h58,8'h93,8'hcf,8'hf4,8'hff,8'hfa,8'hc4,8'h76,8'h98,8'hff,8'hbc,8'h53,8'haa,8'hfb,8'hff,8'he7,8'h76,8'h2a,8'h00,8'h27,8'h27,8'h27,8'h27,8'h27,8'h42,8'he4,8'hee,8'h4f,8'h06,8'h11,8'h3f,8'h97,8'heb,8'hff,8'hff,8'he5,8'h73,8'h2b,8'h25,8'h00,8'h25,8'h59,8'hea,8'hfa,8'h98,8'h3c,8'h2f,8'h48,8'h6c,8'h8f,8'hbb,8'he3,8'hfa,8'hff,8'hfc,8'hec,8'hb0,8'h61,8'h75,8'hee,8'hc2,8'h2c,8'h42,8'hb9,8'hff,8'hfb,8'hb1,8'h40,8'h25,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h72,8'hf0,8'hff,8'hfd,8'hf1,8'he0,8'hb2,8'h92,8'h7b,8'h7f,8'hbe,8'hf5,8'hfc,8'hff,8'hff,8'hff,8'hff,8'hff,8'hf3,8'h7b,8'h0f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h28,8'hb3,8'hff,8'hff,8'hff,8'hff,8'hb6,8'h46,8'h29,8'h31,8'h51,8'h82,8'hbc,8'hec,8'hff,8'hff,8'hfc,8'hde,8'h94,8'h61,8'haf,8'hfb,8'hf8,8'hb4,8'h8c,8'hc7,8'hfb,8'hfa,8'hc5,8'h4c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h25,8'h62,8'he5,8'hff,8'hf5,8'h7a,8'h24,8'h1d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1f,8'h2b,8'h6d,8'hc5,8'hfb,8'hff,8'hff,8'hff,8'hff,8'hd5,8'h31,8'h01,8'h00,8'h00,8'h00,8'h00,8'h16,8'h38,8'h7e,8'hd3,8'hff,8'hff,8'hff,8'hf0,8'hb6,8'h59,8'h30,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h29,8'h8a,8'hf4,8'hff,8'hf0,8'hb5,8'h8f,8'h99,8'haf,8'hd1,8'hef,8'hff,8'hff,8'hf7,8'hdd,8'h87,8'h3d,8'h28,8'h67,8'hf7,8'hfd,8'he9,8'hff,8'hff,8'hcd,8'h66,8'h2c,8'h25,8'h00,8'h27,8'h27,8'h27,8'h27,8'h27,8'h41,8'hdb,8'hff,8'h9a,8'h42,8'h6f,8'hcb,8'hfb,8'hff,8'hfc,8'hd0,8'h6d,8'h2b,8'h26,8'h00,8'h00,8'h25,8'h32,8'h9b,8'hfb,8'hff,8'he4,8'hde,8'hea,8'hfb,8'hff,8'hff,8'hff,8'hef,8'hc8,8'h8f,8'h5e,8'h35,8'h24,8'h4a,8'hd8,8'hf9,8'hbc,8'hd5,8'hff,8'hf3,8'ha7,8'h45,8'h26,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h3c,8'hc0,8'hf6,8'hd9,8'ha3,8'h73,8'h4c,8'h34,8'h2d,8'h28,8'h37,8'ha4,8'hf8,8'hff,8'he7,8'hf8,8'hff,8'hf9,8'hf8,8'hff,8'he3,8'h4a,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h73,8'hfe,8'hff,8'hff,8'hff,8'hff,8'he9,8'hd4,8'hda,8'hef,8'hfe,8'hff,8'hfe,8'hf0,8'hdf,8'ha6,8'h55,8'h2d,8'h27,8'h6b,8'he3,8'hff,8'hff,8'hff,8'hff,8'hfd,8'hc3,8'h54,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h25,8'h35,8'hb0,8'hff,8'hff,8'he4,8'h70,8'h24,8'h0c,8'h1d,8'h17,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h36,8'h6d,8'hba,8'hf5,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hff,8'ha1,8'h13,8'h0b,8'h00,8'h00,8'h1a,8'h3e,8'h74,8'hcd,8'hf9,8'hff,8'hff,8'hf5,8'hc5,8'h77,8'h35,8'h00,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h40,8'hbe,8'hfe,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hf0,8'hdc,8'hb0,8'h73,8'h45,8'h2b,8'h25,8'h00,8'h61,8'he7,8'hff,8'hff,8'hfe,8'hbd,8'h52,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h27,8'h2c,8'h91,8'hff,8'hf5,8'he0,8'hf4,8'hff,8'hff,8'he2,8'h90,8'h4c,8'h28,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h40,8'hb2,8'hf9,8'hff,8'hff,8'hf3,8'he8,8'hdc,8'hc4,8'ha0,8'h65,8'h3b,8'h29,8'h00,8'h26,8'h26,8'h34,8'hb3,8'hfe,8'hff,8'hff,8'hee,8'h93,8'h38,8'h27,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h65,8'hc3,8'h91,8'h4b,8'h2c,8'h27,8'h00,8'h25,8'h25,8'h2c,8'h7c,8'he6,8'hff,8'hd5,8'h8a,8'hed,8'hff,8'hf3,8'hf1,8'hf5,8'hff,8'ha7,8'h21,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h44,8'heb,8'hff,8'hff,8'hdd,8'hd3,8'hf3,8'hff,8'hff,8'hfe,8'hf5,8'he4,8'hb6,8'h71,8'h48,8'h2e,8'h00,8'h25,8'h00,8'h2d,8'h8a,8'he6,8'hfd,8'hff,8'hf2,8'hb7,8'h4f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h66,8'he4,8'hff,8'hff,8'he7,8'h83,8'h3a,8'h20,8'h15,8'h07,8'h0d,8'h0b,8'h00,8'h00,8'h00,8'h0f,8'h22,8'h2b,8'h48,8'h7e,8'hc5,8'hf3,8'hff,8'hff,8'hff,8'hfe,8'hf2,8'hf2,8'hfe,8'hf9,8'h69,8'h09,8'h0a,8'h16,8'h31,8'h73,8'hc8,8'hf6,8'hff,8'hff,8'hf6,8'hd3,8'h8e,8'h43,8'h28,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h55,8'had,8'hc3,8'hd9,8'he4,8'hde,8'hca,8'hbe,8'h82,8'h53,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2f,8'h73,8'hbf,8'hc9,8'ha6,8'h41,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h26,8'h4e,8'hda,8'hff,8'hff,8'hff,8'hff,8'hd3,8'h6b,8'h2a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h4b,8'h8f,8'hb2,8'ha0,8'h74,8'h5c,8'h4e,8'h36,8'h2c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h29,8'h82,8'he8,8'hf7,8'he4,8'h90,8'h39,8'h27,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h4f,8'h54,8'h2c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2a,8'h6c,8'he1,8'hff,8'he9,8'h6b,8'h94,8'hff,8'hfe,8'he6,8'h9d,8'hcf,8'hff,8'he4,8'h3c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h32,8'he2,8'hff,8'hfa,8'h87,8'h4b,8'h84,8'hb5,8'hbb,8'hb5,8'h8a,8'h5d,8'h39,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h35,8'h6f,8'ha8,8'hb2,8'h84,8'h40,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h2e,8'h7b,8'hde,8'hfd,8'hff,8'hf9,8'hd4,8'h8f,8'h5e,8'h43,8'h40,8'h44,8'h46,8'h43,8'h44,8'h59,8'h81,8'hb3,8'hdf,8'hf8,8'hff,8'hff,8'hff,8'hf5,8'hd6,8'haa,8'h7b,8'hba,8'hff,8'he4,8'h3b,8'h22,8'h3e,8'h67,8'hc0,8'hf3,8'hff,8'hff,8'hec,8'hcc,8'h99,8'h56,8'h2e,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h34,8'h3e,8'h4d,8'h5b,8'h54,8'h43,8'h3a,8'h2a,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h28,8'h3a,8'h40,8'h36,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h26,8'h2a,8'h6d,8'hc6,8'hd4,8'hd1,8'ha1,8'h4f,8'h29,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h2c,8'h35,8'h2e,8'h00,8'h24,8'h25,8'h25,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3b,8'h6d,8'h83,8'h5f,8'h33,8'h25,8'h00,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h29,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h28,8'h62,8'hd4,8'hff,8'hed,8'h73,8'h45,8'hdf,8'hff,8'hf4,8'ha3,8'h39,8'h81,8'hf1,8'hfd,8'h71,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h34,8'he3,8'hff,8'hf4,8'h6e,8'h25,8'h2a,8'h36,8'h39,8'h38,8'h2c,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h28,8'h34,8'h36,8'h2a,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h25,8'h2c,8'h53,8'ha1,8'hec,8'hfe,8'hff,8'hff,8'hf3,8'he7,8'he5,8'he5,8'he7,8'he7,8'he7,8'hf0,8'hfd,8'hff,8'hff,8'hff,8'hfb,8'hf2,8'hce,8'h80,8'h44,8'h2f,8'h3a,8'hba,8'hff,8'hc1,8'h59,8'h97,8'hd9,8'hf3,8'hff,8'hff,8'hea,8'hba,8'h65,8'h3e,8'h2d,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h25,8'h24,8'h25,8'h25,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2a,8'h38,8'h3d,8'h3c,8'h2f,8'h25,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h27,8'h29,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h2c,8'h6b,8'hd6,8'hff,8'hef,8'h73,8'h21,8'h93,8'hff,8'hff,8'hd5,8'h51,8'h23,8'h54,8'hda,8'hff,8'ha3,8'h17,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h45,8'heb,8'hff,8'hf1,8'h5c,8'h00,8'h25,8'h25,8'h25,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h31,8'h7b,8'hd7,8'hf7,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hff,8'hfe,8'hed,8'hbd,8'h83,8'h48,8'h2a,8'h25,8'h24,8'h4e,8'hdd,8'hff,8'heb,8'he2,8'hff,8'hff,8'hff,8'hf6,8'hc6,8'h70,8'h36,8'h27,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h27,8'h67,8'hd6,8'hff,8'hf8,8'h7f,8'h18,8'h43,8'he2,8'hff,8'hf9,8'ha0,8'h2e,8'h22,8'h5c,8'hdc,8'hff,8'hbd,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h6c,8'hfd,8'hff,8'hd2,8'h42,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2c,8'h5d,8'h95,8'had,8'hbf,8'hd5,8'he4,8'hf2,8'hf3,8'hf0,8'he8,8'hdb,8'hc6,8'hb2,8'ha7,8'h75,8'h3b,8'h27,8'h00,8'h00,8'h00,8'h00,8'h6d,8'hf3,8'hff,8'hff,8'hff,8'hfe,8'hdb,8'hb2,8'h83,8'h45,8'h28,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2e,8'h65,8'hcf,8'hf9,8'he6,8'h84,8'h21,8'h27,8'h9d,8'hfd,8'hfc,8'hd6,8'h58,8'h3f,8'h73,8'hb8,8'hf7,8'hed,8'h72,8'h0b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1b,8'h9e,8'hff,8'hff,8'h88,8'h2a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h2c,8'h31,8'h3d,8'h4a,8'h5a,8'h6f,8'h76,8'h71,8'h61,8'h4d,8'h41,8'h33,8'h2e,8'h27,8'h25,8'h00,8'h00,8'h00,8'h00,8'h2c,8'h96,8'hff,8'hff,8'hf9,8'he7,8'ha3,8'h55,8'h33,8'h28,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h29,8'h6f,8'hda,8'hff,8'hec,8'h6f,8'h14,8'h06,8'h59,8'he9,8'hff,8'hf4,8'h9d,8'h4a,8'hac,8'hf1,8'hff,8'he8,8'h70,8'h18,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2f,8'hd2,8'hff,8'he8,8'h58,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h25,8'h25,8'h24,8'h25,8'h00,8'h27,8'h00,8'h25,8'h24,8'h25,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3c,8'hc4,8'hf5,8'he5,8'hb1,8'h62,8'h32,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h28,8'h51,8'hc9,8'hfe,8'hed,8'h7b,8'h1b,8'h00,8'h21,8'ha2,8'hff,8'hfd,8'hf8,8'hcd,8'hc2,8'hf9,8'hff,8'hd4,8'h61,8'h12,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h18,8'h6f,8'hf7,8'hff,8'hb2,8'h35,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h51,8'ha4,8'h7a,8'h52,8'h32,8'h27,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h2f,8'h75,8'hd1,8'hfd,8'hda,8'h65,8'h1d,8'h00,8'h05,8'h65,8'hf1,8'hff,8'hf5,8'hf8,8'hfb,8'hff,8'he7,8'h8d,8'h42,8'h08,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h41,8'hcd,8'hff,8'hef,8'h6d,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3d,8'h3d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h38,8'h87,8'he9,8'hff,8'hd2,8'h4f,8'h01,8'h00,8'h00,8'h31,8'hc5,8'hff,8'hf6,8'hf6,8'hff,8'hff,8'hcd,8'h58,8'h13,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h99,8'hff,8'hff,8'hb3,8'h39,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3f,8'h9c,8'hed,8'hfa,8'hcf,8'h53,8'h0b,8'h00,8'h00,8'h0f,8'h7a,8'hf9,8'hfd,8'hfa,8'hfe,8'hed,8'ha8,8'h39,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h72,8'hf1,8'hff,8'he3,8'h5f,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h29,8'h59,8'hbd,8'hf5,8'hfb,8'ha2,8'h3c,8'h06,8'h00,8'h00,8'h00,8'h52,8'hdf,8'hff,8'hff,8'hf0,8'ha7,8'h4a,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h8b,8'hed,8'hff,8'hea,8'h72,8'h2b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2e,8'h6f,8'hd6,8'hff,8'hfa,8'h9d,8'h27,8'h00,8'h00,8'h00,8'h00,8'h29,8'hb2,8'hff,8'hfe,8'hc9,8'h64,8'h22,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h28,8'h8a,8'hf5,8'hff,8'hf3,8'h8a,8'h2d,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h5e,8'hdb,8'hfb,8'he0,8'h8a,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h62,8'hd2,8'hc7,8'h84,8'h35,8'h02,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0d,8'h3b,8'h9a,8'hf2,8'hff,8'hec,8'h96,8'h39,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h6f,8'hef,8'hf7,8'h76,8'h19,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h39,8'h46,8'h28,8'h18,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h22,8'h47,8'hbf,8'hfd,8'hff,8'he7,8'h80,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h64,8'hec,8'hf8,8'h62,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h05,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1d,8'h53,8'hca,8'hff,8'hff,8'he5,8'h76,8'h2e,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h64,8'hec,8'hfe,8'h71,8'h08,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2c,8'h7a,8'he1,8'hff,8'hfe,8'hca,8'h6e,8'h2c,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h60,8'he7,8'hff,8'h82,8'h1a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h34,8'h9c,8'hf5,8'hff,8'hfe,8'hc2,8'h4e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h4d,8'hda,8'hff,8'h92,8'h21,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0c,8'h3e,8'hb1,8'hff,8'hff,8'hf7,8'hbd,8'h4e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h3a,8'hcb,8'hff,8'hae,8'h22,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h6d,8'hd1,8'hff,8'hff,8'hea,8'h92,8'h3f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h38,8'hca,8'hff,8'hb3,8'h1f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h2d,8'h90,8'hf0,8'hff,8'hff,8'hde,8'h70,8'h2f,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h37,8'hc7,8'hff,8'hba,8'h23,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h12,8'h3f,8'hae,8'hfb,8'hff,8'hfa,8'hcc,8'h6b,8'h2b,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h32,8'hb9,8'hff,8'hc3,8'h2a,8'h02,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h18,8'h58,8'hc6,8'hff,8'hff,8'hf4,8'hb2,8'h4c,8'h29,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2c,8'ha2,8'hff,8'hd3,8'h36,8'h03,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h02,8'h25,8'h75,8'he2,8'hff,8'hff,8'hf3,8'hac,8'h42,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h8e,8'hfc,8'hdc,8'h3e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h21,8'h3f,8'h9a,8'hf3,8'hff,8'hf9,8'hdb,8'h8f,8'h3d,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8d,8'hf9,8'he2,8'h42,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0d,8'h2e,8'h7b,8'hd2,8'hfc,8'hff,8'hf0,8'hac,8'h53,8'h2e,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8f,8'hfc,8'he5,8'h42,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'h00,8'h0b,8'h40,8'ha9,8'hf6,8'hff,8'hfe,8'he3,8'h89,8'h3b,8'h25,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8f,8'hfd,8'he5,8'h43,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h14,8'h2f,8'h6f,8'hd4,8'hff,8'hff,8'hf1,8'hc0,8'h65,8'h2e,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8e,8'hfb,8'he1,8'h44,8'h05,8'h08,8'h01,8'h05,8'h01,8'h1c,8'h5f,8'hc8,8'hf9,8'hfe,8'hfb,8'hdb,8'h83,8'h39,8'h27,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8e,8'hfb,8'he3,8'h43,8'h10,8'h0e,8'h10,8'h1a,8'h36,8'h8b,8'he6,8'hff,8'hfc,8'hf4,8'hc2,8'h64,8'h2b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8f,8'hfb,8'he1,8'h44,8'h19,8'h12,8'h39,8'h7b,8'hc6,8'hf6,8'hfd,8'hf5,8'hd6,8'h93,8'h47,8'h27,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8f,8'hf9,8'hd7,8'h3c,8'h1a,8'h52,8'hc2,8'hf9,8'hff,8'hfc,8'he6,8'ha2,8'h4e,8'h2d,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8f,8'hfb,8'hdc,8'h61,8'h83,8'he5,8'hfe,8'hfa,8'he9,8'hc4,8'h70,8'h32,8'h00,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h8f,8'hf8,8'hf8,8'he0,8'hf0,8'hfb,8'hee,8'hc3,8'h7c,8'h43,8'h28,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h92,8'hf8,8'hff,8'hff,8'hfc,8'hed,8'hab,8'h4d,8'h28,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2d,8'ha6,8'hfa,8'hfa,8'hec,8'hd6,8'h87,8'h3c,8'h00,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h32,8'hb8,8'hf4,8'hc6,8'h72,8'h45,8'h2b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h34,8'hb5,8'haa,8'h4b,8'h28,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2a,8'h4d,8'h3c,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}};

parameter bit [7:0] SpriteTableG[111:0][226:0] = '{'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h27,8'h27,8'h26,8'h26,8'h23,8'h24,8'h23,8'h22,8'h1c,8'h1a,8'h18,8'h14,8'h19,8'h19,8'h17,8'h19,8'h19,8'h19,8'h19,8'h16,8'h19,8'h1c,8'h1c,8'h18,8'h19,8'h1b,8'h20,8'h22,8'h23,8'h22,8'h21,8'h24,8'h26,8'h26,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h26,8'h25,8'h23,8'h23,8'h24,8'h21,8'h12,8'h09,8'h08,8'h0c,8'h0f,8'h16,8'h17,8'h21,8'h26,8'h2f,8'h35,8'h37,8'h3a,8'h3a,8'h3a,8'h38,8'h37,8'h37,8'h39,8'h3f,8'h3e,8'h3a,8'h39,8'h3e,8'h39,8'h36,8'h2f,8'h29,8'h22,8'h23,8'h1d,8'h1a,8'h24,8'h25,8'h23,8'h24,8'h24,8'h25,8'h26,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h00,8'h27,8'h26,8'h25,8'h24,8'h22,8'h18,8'h06,8'h00,8'h00,8'h00,8'h1b,8'h2f,8'h3a,8'h45,8'h54,8'h5c,8'h62,8'h6b,8'h6c,8'h6c,8'h69,8'h64,8'h65,8'h62,8'h59,8'h53,8'h56,8'h55,8'h55,8'h50,8'h55,8'h55,8'h55,8'h5a,8'h5c,8'h60,8'h6a,8'h69,8'h67,8'h69,8'h6f,8'h70,8'h6b,8'h65,8'h5c,8'h55,8'h49,8'h39,8'h29,8'h13,8'h0d,8'h0c,8'h12,8'h21,8'h23,8'h24,8'h25,8'h26,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h27,8'h25,8'h23,8'h21,8'h19,8'h00,8'h00,8'h00,8'h15,8'h2d,8'h40,8'h48,8'h57,8'h63,8'h69,8'h6b,8'h66,8'h61,8'h60,8'h54,8'h4b,8'h4e,8'h4a,8'h44,8'h46,8'h49,8'h4f,8'h54,8'h55,8'h59,8'h5b,8'h59,8'h5c,8'h5d,8'h61,8'h5d,8'h58,8'h56,8'h58,8'h54,8'h4e,8'h47,8'h46,8'h47,8'h49,8'h4b,8'h48,8'h4e,8'h5d,8'h62,8'h64,8'h6d,8'h6b,8'h6b,8'h65,8'h53,8'h43,8'h2f,8'h24,8'h0d,8'h0b,8'h0e,8'h1b,8'h22,8'h24,8'h25,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h26,8'h23,8'h23,8'h1a,8'h00,8'h00,8'h00,8'h21,8'h3e,8'h53,8'h63,8'h6a,8'h66,8'h69,8'h62,8'h54,8'h4b,8'h46,8'h48,8'h4d,8'h59,8'h65,8'h70,8'h7a,8'h88,8'h93,8'h96,8'ha2,8'had,8'hae,8'hb4,8'hb5,8'hba,8'hb7,8'hb8,8'hbb,8'hbd,8'hbf,8'hbd,8'hba,8'hb7,8'hbb,8'hb4,8'haf,8'ha7,8'ha4,8'h9d,8'h99,8'h90,8'h81,8'h75,8'h68,8'h5d,8'h4e,8'h4c,8'h4b,8'h51,8'h56,8'h5d,8'h64,8'h68,8'h6b,8'h66,8'h5b,8'h42,8'h2a,8'h12,8'h00,8'h0f,8'h20,8'h24,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h00,8'h27,8'h26,8'h25,8'h23,8'h10,8'h00,8'h00,8'h20,8'h3b,8'h52,8'h65,8'h70,8'h6f,8'h61,8'h53,8'h48,8'h43,8'h4d,8'h5e,8'h6e,8'h81,8'h93,8'ha3,8'haf,8'hbb,8'hbd,8'hc0,8'hc4,8'hc5,8'hc8,8'hc3,8'hc2,8'hc1,8'hb8,8'hb6,8'hb1,8'hb0,8'ha8,8'ha5,8'ha5,8'ha5,8'ha5,8'ha2,8'ha0,8'ha1,8'ha3,8'ha7,8'had,8'hae,8'hb0,8'hb6,8'hbd,8'hc2,8'hc3,8'hc2,8'hbd,8'hb7,8'haf,8'ha6,8'h99,8'h86,8'h75,8'h67,8'h58,8'h4b,8'h4b,8'h52,8'h5f,8'h67,8'h6e,8'h6b,8'h5b,8'h45,8'h25,8'h09,8'h17,8'h21,8'h25,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h27,8'h25,8'h24,8'h20,8'h06,8'h00,8'h00,8'h24,8'h43,8'h5c,8'h73,8'h74,8'h60,8'h4b,8'h49,8'h4f,8'h5c,8'h71,8'h89,8'ha4,8'had,8'hb9,8'hc5,8'hc5,8'hc6,8'hc4,8'hc7,8'hc0,8'hb2,8'had,8'ha2,8'h94,8'h85,8'h79,8'h6e,8'h65,8'h58,8'h4d,8'h48,8'h48,8'h45,8'h42,8'h42,8'h41,8'h42,8'h40,8'h3f,8'h40,8'h3f,8'h44,8'h47,8'h47,8'h4b,8'h52,8'h5b,8'h65,8'h74,8'h80,8'h89,8'h98,8'ha6,8'had,8'hb4,8'hb8,8'hb7,8'hb5,8'hb0,8'ha4,8'h91,8'h78,8'h5f,8'h4d,8'h45,8'h4a,8'h5c,8'h6e,8'h73,8'h61,8'h47,8'h2c,8'h12,8'h11,8'h22,8'h23,8'h26,8'h26,8'h26,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h26,8'h24,8'h1c,8'h10,8'h00,8'h03,8'h2f,8'h4a,8'h4b,8'h4d,8'h54,8'h62,8'h67,8'h6e,8'h75,8'h73,8'h7b,8'h9a,8'hb1,8'hc2,8'hc8,8'hc7,8'hc4,8'hb6,8'ha3,8'h88,8'h72,8'h6e,8'h71,8'h70,8'h66,8'h5f,8'h57,8'h54,8'h55,8'h53,8'h4f,8'h49,8'h48,8'h47,8'h46,8'h44,8'h47,8'h4a,8'h4e,8'h55,8'h51,8'h50,8'h54,8'h51,8'h4e,8'h4e,8'h50,8'h4c,8'h4a,8'h48,8'h49,8'h47,8'h48,8'h4d,8'h50,8'h59,8'h57,8'h5a,8'h59,8'h63,8'h6c,8'h73,8'h73,8'h70,8'h7c,8'h8e,8'ha5,8'hae,8'had,8'h9f,8'h84,8'h74,8'h70,8'h66,8'h64,8'h63,8'h53,8'h51,8'h4e,8'h4a,8'h36,8'h24,8'h21,8'h26,8'h24,8'h26,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h25,8'h1c,8'h00,8'h00,8'h00,8'h29,8'h4d,8'h63,8'h69,8'h61,8'h50,8'h4e,8'h59,8'h7b,8'ha2,8'hbb,8'hca,8'hcc,8'hcc,8'hc5,8'hbe,8'hac,8'h8f,8'h72,8'h5f,8'h4a,8'h3d,8'h36,8'h39,8'h41,8'h4e,8'h55,8'h5e,8'h65,8'h66,8'h60,8'h5b,8'h58,8'h4f,8'h47,8'h40,8'h31,8'h2a,8'h26,8'h21,8'h13,8'h0e,8'h05,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1a,8'h22,8'h29,8'h30,8'h37,8'h40,8'h45,8'h4e,8'h50,8'h55,8'h53,8'h5a,8'h57,8'h51,8'h52,8'h46,8'h42,8'h41,8'h43,8'h56,8'h6a,8'h81,8'h9b,8'hb6,8'hc0,8'hb7,8'ha0,8'h79,8'h58,8'h46,8'h4a,8'h60,8'h65,8'h2f,8'h25,8'h5b,8'h2b,8'h0b,8'h21,8'h25,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h23,8'h20,8'h14,8'h00,8'h0a,8'h3f,8'h5e,8'h6a,8'h65,8'h55,8'h50,8'h65,8'h85,8'ha7,8'hbe,8'hcb,8'hcc,8'hc3,8'hbf,8'haf,8'h93,8'h71,8'h5f,8'h46,8'h3a,8'h3d,8'h47,8'h4c,8'h59,8'h63,8'h65,8'h63,8'h54,8'h45,8'h35,8'h29,8'h1c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h23,8'h0e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h11,8'h26,8'h33,8'h43,8'h4b,8'h57,8'h5a,8'h52,8'h52,8'h49,8'h40,8'h47,8'h50,8'h6a,8'h87,8'h9d,8'hb6,8'hb5,8'h9c,8'h7d,8'h4a,8'h28,8'h22,8'h3f,8'h84,8'h73,8'h46,8'h22,8'h22,8'h25,8'h25,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h26,8'h24,8'h26,8'h26,8'h24,8'h24,8'h24,8'h25,8'h26,8'h27,8'h27,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h26,8'h24,8'h20,8'h08,8'h00,8'h2a,8'h55,8'h61,8'h4e,8'h46,8'h5a,8'h6e,8'h8b,8'h9b,8'haa,8'hc4,8'hcc,8'hc6,8'hb8,8'h9b,8'h74,8'h53,8'h4c,8'h52,8'h50,8'h56,8'h66,8'h61,8'h56,8'h51,8'h42,8'h2d,8'h2b,8'h24,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'h0c,8'h11,8'h18,8'h16,8'h1c,8'h1c,8'h21,8'h22,8'h25,8'h22,8'h36,8'h29,8'h28,8'h29,8'h2b,8'h33,8'h31,8'h24,8'h3b,8'h37,8'h25,8'h26,8'h24,8'h2b,8'h1c,8'h25,8'h26,8'h16,8'h11,8'h18,8'h19,8'h14,8'h11,8'h07,8'h00,8'h00,8'h00,8'h00,8'h00,8'h19,8'h28,8'h30,8'h31,8'h40,8'h4b,8'h60,8'h68,8'h63,8'h61,8'h57,8'h62,8'h78,8'h55,8'h2f,8'h64,8'h9d,8'h92,8'h6d,8'h52,8'h59,8'h66,8'h59,8'h37,8'h25,8'h21,8'h24,8'h26,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h00,8'h25,8'h23,8'h21,8'h20,8'h20,8'h2b,8'h38,8'h46,8'h51,8'h5a,8'h5e,8'h5d,8'h56,8'h4f,8'h34,8'h22,8'h26,8'h27,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h26,8'h22,8'h03,8'h00,8'h00,8'h32,8'h5e,8'h69,8'h5b,8'h45,8'h4c,8'h77,8'ha6,8'hc2,8'hcd,8'hcd,8'hc3,8'hb2,8'h91,8'h6b,8'h4c,8'h34,8'h36,8'h4c,8'h5f,8'h6c,8'h68,8'h58,8'h42,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0c,8'h14,8'h15,8'h1b,8'h21,8'h21,8'h22,8'h20,8'h20,8'h21,8'h21,8'h25,8'h30,8'h39,8'h43,8'h2c,8'h28,8'h2b,8'h48,8'h4b,8'h22,8'h50,8'h54,8'h38,8'h33,8'h4d,8'h44,8'h25,8'h22,8'h25,8'h2f,8'h43,8'h42,8'h2c,8'h20,8'h20,8'h20,8'h20,8'h21,8'h22,8'h22,8'h23,8'h24,8'h24,8'h13,8'h0c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2d,8'h48,8'h58,8'h56,8'h3b,8'h31,8'h4e,8'h38,8'h72,8'hb5,8'hc0,8'hba,8'h92,8'h66,8'h5a,8'h68,8'h73,8'h65,8'h41,8'h22,8'h1f,8'h23,8'h25,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h25,8'h23,8'h20,8'h14,8'h21,8'h30,8'h4e,8'h68,8'h7b,8'h83,8'h7e,8'h78,8'h78,8'h78,8'h78,8'h83,8'h90,8'h89,8'h47,8'h1e,8'h26,8'h27},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h26,8'h24,8'h13,8'h06,8'h1e,8'h31,8'h4c,8'h67,8'h67,8'h5a,8'h5e,8'h86,8'hb4,8'hc5,8'hc2,8'hbb,8'ha3,8'h8f,8'h78,8'h5e,8'h45,8'h40,8'h4a,8'h54,8'h63,8'h63,8'h4f,8'h2c,8'h00,8'h00,8'h00,8'h00,8'h08,8'h1a,8'h25,8'h22,8'h1d,8'h18,8'h1d,8'h20,8'h20,8'h1b,8'h1a,8'h21,8'h21,8'h22,8'h23,8'h23,8'h24,8'h24,8'h24,8'h27,8'h34,8'h40,8'h3c,8'h35,8'h30,8'h32,8'h30,8'h27,8'h35,8'h3a,8'h4d,8'h3f,8'h46,8'h3e,8'h26,8'h2d,8'h43,8'h7b,8'hae,8'h9c,8'h60,8'h33,8'h28,8'h22,8'h25,8'h31,8'h2c,8'h2b,8'h2c,8'h35,8'h30,8'h21,8'h24,8'h23,8'h20,8'h2b,8'h2d,8'h23,8'h00,8'h00,8'h00,8'h00,8'h24,8'h4b,8'h69,8'h4a,8'h3b,8'h40,8'h57,8'h76,8'h92,8'ha5,8'ha6,8'h99,8'h77,8'h64,8'h7d,8'h7a,8'h60,8'h47,8'h37,8'h2e,8'h27,8'h26,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h26,8'h25,8'h28,8'h2c,8'h36,8'h48,8'h5f,8'h74,8'h79,8'h6e,8'h64,8'h5d,8'h53,8'h4d,8'h48,8'h47,8'h47,8'h4d,8'h53,8'h77,8'h83,8'h29,8'h20,8'h26},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h25,8'h20,8'h00,8'h04,8'h39,8'h5e,8'h61,8'h46,8'h4e,8'h79,8'h9a,8'haf,8'hbc,8'hc9,8'hc7,8'hac,8'h79,8'h51,8'h3e,8'h48,8'h5b,8'h69,8'h60,8'h4c,8'h37,8'h21,8'h00,8'h00,8'h00,8'h00,8'h06,8'h0f,8'h29,8'h50,8'h35,8'h27,8'h32,8'h27,8'h11,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1e,8'h21,8'h21,8'h23,8'h24,8'h24,8'h24,8'h24,8'h23,8'h26,8'h29,8'h3b,8'h32,8'h33,8'h28,8'h2c,8'h33,8'h41,8'h26,8'h2d,8'h40,8'h45,8'h32,8'h2b,8'h38,8'h4b,8'h89,8'he7,8'hc1,8'h5c,8'h43,8'h31,8'h25,8'h25,8'h3e,8'h4a,8'h2e,8'h23,8'h26,8'h25,8'h23,8'h28,8'h23,8'h24,8'h3f,8'h49,8'h50,8'h34,8'h2b,8'h2a,8'h0d,8'h34,8'h83,8'h57,8'h25,8'h02,8'h26,8'h43,8'h5e,8'h61,8'h5a,8'h54,8'h69,8'h93,8'haa,8'hac,8'h8f,8'h6a,8'h5e,8'h6b,8'h72,8'h50,8'h28,8'h22,8'h25,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h25,8'h24,8'h2c,8'h47,8'h67,8'h6d,8'h59,8'h48,8'h45,8'h5a,8'h70,8'h7f,8'h91,8'ha0,8'ha8,8'hac,8'haf,8'hb1,8'hb1,8'haf,8'h90,8'h44,8'h7a,8'h51,8'h0c,8'h26},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h25,8'h1a,8'h00,8'h00,8'h38,8'h62,8'h67,8'h48,8'h4c,8'h75,8'ha7,8'hc3,8'hca,8'hce,8'hbd,8'ha1,8'h70,8'h45,8'h39,8'h4b,8'h61,8'h69,8'h61,8'h3d,8'h0b,8'h00,8'h00,8'h00,8'h26,8'h25,8'h24,8'h1f,8'h21,8'h1e,8'h25,8'h3b,8'h29,8'h22,8'h20,8'h00,8'h00,8'h00,8'h00,8'h1d,8'h1a,8'h00,8'h00,8'h0e,8'h21,8'h23,8'h23,8'h23,8'h24,8'h24,8'h24,8'h24,8'h27,8'h28,8'h24,8'h23,8'h22,8'h24,8'h24,8'h24,8'h2b,8'h24,8'h2b,8'h2d,8'h34,8'h2d,8'h22,8'h23,8'h28,8'h4d,8'h95,8'h85,8'h50,8'h24,8'h21,8'h22,8'h24,8'h28,8'h33,8'h28,8'h21,8'h21,8'h25,8'h45,8'h34,8'h3a,8'h49,8'h31,8'h2f,8'h38,8'h2d,8'h48,8'h3c,8'h2d,8'h88,8'h7b,8'h40,8'h22,8'h00,8'h00,8'h00,8'h03,8'h32,8'h52,8'h61,8'h53,8'h46,8'h53,8'h82,8'hac,8'hb0,8'h8f,8'h60,8'h5c,8'h74,8'h70,8'h43,8'h23,8'h23,8'h25,8'h26,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h25,8'h23,8'h2a,8'h4e,8'h72,8'h70,8'h52,8'h3e,8'h4a,8'h6e,8'h95,8'ha1,8'ha2,8'h93,8'h7d,8'h6d,8'h92,8'hc5,8'hd0,8'hce,8'hce,8'hcf,8'hb6,8'h42,8'h6c,8'h53,8'h17,8'h27},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h25,8'h21,8'h0b,8'h24,8'h3c,8'h4e,8'h68,8'h69,8'h61,8'h73,8'haf,8'hca,8'hc7,8'hbc,8'h9c,8'h82,8'h65,8'h4e,8'h43,8'h4f,8'h60,8'h5c,8'h4a,8'h25,8'h00,8'h00,8'h00,8'h1c,8'h2e,8'h33,8'h52,8'h40,8'h28,8'h22,8'h22,8'h22,8'h21,8'h1a,8'h11,8'h00,8'h00,8'h00,8'h23,8'h24,8'h35,8'h55,8'h62,8'h45,8'h00,8'h00,8'h1e,8'h21,8'h24,8'h26,8'h23,8'h23,8'h24,8'h24,8'h23,8'h23,8'h22,8'h21,8'h22,8'h23,8'h22,8'h21,8'h21,8'h21,8'h25,8'h23,8'h21,8'h23,8'h22,8'h23,8'h26,8'h29,8'h4c,8'h4b,8'h3f,8'h26,8'h23,8'h22,8'h24,8'h31,8'h32,8'h29,8'h23,8'h24,8'h28,8'h4b,8'h3a,8'h45,8'h4b,8'h33,8'h30,8'h36,8'h2d,8'h27,8'h45,8'h8c,8'h7e,8'h39,8'h3a,8'h24,8'h22,8'h22,8'h16,8'h00,8'h00,8'h00,8'h00,8'h3f,8'h53,8'h45,8'h43,8'h60,8'h7b,8'h8e,8'h9b,8'h86,8'h6d,8'h77,8'h73,8'h57,8'h45,8'h32,8'h21,8'h24,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h25,8'h23,8'h2a,8'h41,8'h4f,8'h64,8'h6e,8'h68,8'h60,8'h66,8'h8a,8'h9a,8'h8e,8'h89,8'h6f,8'h5d,8'h4b,8'h45,8'h3e,8'h42,8'ha8,8'hd0,8'hca,8'hcb,8'hc8,8'h8d,8'h43,8'h71,8'h30,8'h16,8'h26},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h27,8'h26,8'h24,8'h25,8'h26,8'h24,8'h23,8'h26,8'h25,8'h26,8'h00,8'h27,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h22,8'h0c,8'h23,8'h4f,8'h67,8'h57,8'h4a,8'h67,8'ha2,8'hc2,8'hcb,8'hc8,8'hb7,8'h8e,8'h60,8'h3d,8'h46,8'h60,8'h67,8'h54,8'h3e,8'h00,8'h00,8'h00,8'h00,8'h1a,8'h1a,8'h1f,8'h28,8'h2e,8'h2b,8'h22,8'h25,8'h22,8'h20,8'h22,8'h20,8'h00,8'h00,8'h00,8'h00,8'h2f,8'h42,8'h42,8'h3d,8'h50,8'h4e,8'h38,8'h63,8'h09,8'h00,8'h1f,8'h26,8'h34,8'h4c,8'h33,8'h2b,8'h24,8'h21,8'h21,8'h22,8'h22,8'h21,8'h21,8'h22,8'h22,8'h22,8'h21,8'h21,8'h23,8'h23,8'h23,8'h24,8'h23,8'h24,8'h23,8'h22,8'h34,8'h34,8'h21,8'h2b,8'h38,8'h24,8'h21,8'h30,8'h30,8'h25,8'h24,8'h24,8'h24,8'h2c,8'h41,8'h3e,8'h51,8'h32,8'h44,8'h53,8'h24,8'h45,8'hb4,8'h97,8'h2a,8'h20,8'h25,8'h24,8'h23,8'h24,8'h24,8'h22,8'h21,8'h1f,8'h0d,8'h00,8'h00,8'h00,8'h30,8'h4b,8'h52,8'h4f,8'h54,8'h71,8'h9a,8'ha4,8'h7f,8'h5b,8'h63,8'h6d,8'h4c,8'h25,8'h22,8'h25,8'h00,8'h00,8'h00,8'h27,8'h26,8'h24,8'h25,8'h3c,8'h69,8'h70,8'h53,8'h4d,8'h6c,8'ha4,8'hc4,8'hb0,8'h81,8'h53,8'h4c,8'h60,8'h64,8'h5b,8'h48,8'h45,8'h6b,8'h49,8'h96,8'hd3,8'hce,8'hce,8'hb6,8'h51,8'h61,8'h61,8'h0d,8'h23,8'h27},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h25,8'h23,8'h21,8'h16,8'h0d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h05,8'h17,8'h21,8'h23,8'h25,8'h27,8'h27,8'h26,8'h23,8'h06,8'h05,8'h43,8'h68,8'h5e,8'h49,8'h64,8'h9e,8'hc2,8'hc7,8'hc7,8'hc0,8'h90,8'h59,8'h37,8'h3d,8'h60,8'h68,8'h50,8'h2e,8'h00,8'h00,8'h00,8'h02,8'h1b,8'h21,8'h23,8'h21,8'h24,8'h2b,8'h28,8'h22,8'h20,8'h20,8'h20,8'h20,8'h06,8'h00,8'h00,8'h00,8'h34,8'h4d,8'h42,8'h3a,8'h60,8'h8e,8'hb6,8'h9f,8'h3e,8'h5b,8'h05,8'h00,8'h28,8'h4b,8'h51,8'h46,8'h47,8'h50,8'h31,8'h26,8'h21,8'h22,8'h22,8'h21,8'h21,8'h21,8'h21,8'h21,8'h21,8'h22,8'h23,8'h24,8'h24,8'h24,8'h24,8'h25,8'h23,8'h25,8'h32,8'h2c,8'h24,8'h25,8'h2d,8'h25,8'h21,8'h21,8'h24,8'h24,8'h24,8'h23,8'h25,8'h2c,8'h2c,8'h28,8'h38,8'h2c,8'h30,8'h32,8'h41,8'hb1,8'hc0,8'h45,8'h1e,8'h2a,8'h2b,8'h23,8'h24,8'h24,8'h24,8'h24,8'h26,8'h53,8'h45,8'h22,8'h1e,8'h07,8'h00,8'h00,8'h13,8'h40,8'h53,8'h56,8'h4b,8'h68,8'h9c,8'h9f,8'h71,8'h56,8'h61,8'h68,8'h44,8'h23,8'h22,8'h26,8'h27,8'h25,8'h22,8'h32,8'h5f,8'h6f,8'h5a,8'h4e,8'h71,8'ha3,8'hc6,8'hc9,8'h94,8'h54,8'h4e,8'h62,8'h5f,8'h44,8'h23,8'h00,8'h00,8'h00,8'h53,8'h4b,8'ha7,8'hd5,8'hd0,8'hcd,8'h85,8'h42,8'h7b,8'h2f,8'h19,8'h27,8'h27},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h00,8'h26,8'h24,8'h21,8'h09,8'h00,8'h00,8'h00,8'h24,8'h47,8'h60,8'h65,8'h66,8'h65,8'h67,8'h6a,8'h6d,8'h69,8'h56,8'h32,8'h21,8'h18,8'h07,8'h00,8'h09,8'h4b,8'h5f,8'h52,8'h5f,8'h7c,8'ha1,8'hc5,8'hcd,8'hc8,8'ha9,8'h74,8'h55,8'h4c,8'h57,8'h5a,8'h49,8'h35,8'h19,8'h00,8'h00,8'h16,8'h1f,8'h21,8'h21,8'h23,8'h21,8'h21,8'h23,8'h27,8'h28,8'h22,8'h1e,8'h1d,8'h1f,8'h05,8'h00,8'h00,8'h0e,8'h41,8'h3a,8'h48,8'h67,8'h80,8'h9a,8'hbe,8'hc5,8'hc8,8'ha9,8'h42,8'h57,8'h1f,8'h00,8'h31,8'h35,8'h34,8'h2e,8'h4c,8'h77,8'h37,8'h25,8'h22,8'h22,8'h22,8'h21,8'h21,8'h21,8'h22,8'h22,8'h23,8'h23,8'h24,8'h24,8'h23,8'h23,8'h33,8'h41,8'h3b,8'h29,8'h2f,8'h2b,8'h2f,8'h3c,8'h2a,8'h22,8'h23,8'h24,8'h24,8'h24,8'h24,8'h25,8'h2c,8'h30,8'h2b,8'h25,8'h27,8'h26,8'h27,8'h4e,8'hb2,8'hbf,8'h4b,8'h20,8'h21,8'h39,8'h45,8'h21,8'h23,8'h22,8'h23,8'h28,8'h2b,8'h45,8'h38,8'h28,8'h27,8'h2c,8'h3f,8'h2c,8'h24,8'h00,8'h00,8'h2c,8'h37,8'h4f,8'h6a,8'h6a,8'h75,8'h8a,8'h82,8'h6a,8'h53,8'h55,8'h49,8'h29,8'h23,8'h3f,8'h54,8'h51,8'h55,8'h6e,8'h88,8'hab,8'hc8,8'hc9,8'ha1,8'h69,8'h62,8'h57,8'h47,8'h2f,8'h02,8'h08,8'h1d,8'h21,8'h0c,8'h26,8'h4c,8'h5a,8'hc4,8'hce,8'hca,8'ha4,8'h4c,8'h61,8'h4f,8'h09,8'h25,8'h27,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h26,8'h23,8'h04,8'h00,8'h00,8'h00,8'h29,8'h53,8'h72,8'h85,8'h8a,8'h7e,8'h6c,8'h60,8'h52,8'h4d,8'h4f,8'h60,8'h74,8'h88,8'h8b,8'h74,8'h4d,8'h16,8'h2e,8'h66,8'h67,8'h49,8'h67,8'hab,8'hcc,8'hd2,8'hcc,8'hb4,8'h82,8'h44,8'h36,8'h4f,8'h66,8'h56,8'h27,8'h00,8'h00,8'h00,8'h0e,8'h20,8'h22,8'h24,8'h27,8'h23,8'h22,8'h26,8'h23,8'h2e,8'h28,8'h21,8'h21,8'h18,8'h00,8'h00,8'h00,8'h00,8'h3e,8'h45,8'h3f,8'h50,8'h8b,8'hbb,8'hc8,8'hca,8'hc9,8'hc2,8'hc4,8'ha7,8'h43,8'h55,8'h23,8'h21,8'h43,8'h21,8'h25,8'h26,8'h2a,8'h3a,8'h23,8'h20,8'h23,8'h22,8'h21,8'h21,8'h22,8'h26,8'h27,8'h26,8'h23,8'h21,8'h22,8'h23,8'h22,8'h30,8'h4a,8'h44,8'h39,8'h30,8'h2a,8'h28,8'h27,8'h36,8'h2c,8'h22,8'h24,8'h24,8'h24,8'h24,8'h23,8'h24,8'h2a,8'h37,8'h28,8'h22,8'h22,8'h22,8'h4b,8'hc7,8'hdb,8'h54,8'h17,8'h25,8'h2a,8'h41,8'h57,8'h24,8'h26,8'h24,8'h24,8'h26,8'h25,8'h22,8'h2b,8'h56,8'h4f,8'h47,8'h61,8'h40,8'h41,8'h36,8'h21,8'h00,8'h00,8'h00,8'h3e,8'h56,8'h4c,8'h55,8'h81,8'h9a,8'h76,8'h4d,8'h60,8'h62,8'h57,8'h62,8'h47,8'h48,8'h84,8'hbe,8'hcd,8'hcc,8'hc5,8'h8c,8'h4c,8'h57,8'h5c,8'h25,8'h00,8'h06,8'h20,8'h25,8'h27,8'h26,8'h21,8'h48,8'h46,8'h88,8'hd1,8'hd0,8'hbd,8'h5d,8'h4b,8'h61,8'h04,8'h23,8'h27,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h25,8'h15,8'h00,8'h00,8'h21,8'h45,8'h67,8'h7f,8'h82,8'h76,8'h61,8'h52,8'h5e,8'h6b,8'h7c,8'h8a,8'h8b,8'h82,8'h6e,8'h57,8'h4e,8'h60,8'h76,8'h81,8'h71,8'h65,8'h5b,8'h5e,8'h93,8'hc2,8'hcc,8'hc6,8'hb8,8'h90,8'h60,8'h3f,8'h44,8'h61,8'h55,8'h26,8'h00,8'h00,8'h23,8'h1d,8'h21,8'h22,8'h21,8'h22,8'h26,8'h2c,8'h25,8'h2a,8'h4f,8'h34,8'h26,8'h22,8'h20,8'h14,8'h00,8'h00,8'h00,8'h22,8'h41,8'h34,8'h31,8'h6b,8'hb0,8'hcc,8'hca,8'hc8,8'hc9,8'hc7,8'hc6,8'hc6,8'ha7,8'h44,8'h58,8'h20,8'h03,8'h2b,8'h20,8'h26,8'h28,8'h21,8'h23,8'h22,8'h22,8'h23,8'h21,8'h26,8'h2b,8'h28,8'h3f,8'h3e,8'h32,8'h22,8'h22,8'h24,8'h28,8'h26,8'h2e,8'h2d,8'h2f,8'h3c,8'h38,8'h28,8'h2e,8'h22,8'h24,8'h25,8'h24,8'h24,8'h23,8'h24,8'h25,8'h24,8'h24,8'h25,8'h26,8'h24,8'h22,8'h24,8'h50,8'hc6,8'he8,8'h7d,8'h27,8'h26,8'h3a,8'h5d,8'h8f,8'ha0,8'h61,8'h3b,8'h2e,8'h3b,8'h37,8'h25,8'h22,8'h2c,8'h36,8'h3c,8'h5e,8'h46,8'h4b,8'h58,8'h3d,8'h29,8'h3a,8'h25,8'h08,8'h00,8'h0d,8'h41,8'h4f,8'h48,8'h60,8'h8d,8'h84,8'h5f,8'h58,8'h57,8'h4b,8'h71,8'hae,8'hc9,8'hcb,8'hcc,8'hb7,8'h7d,8'h50,8'h5c,8'h50,8'h13,8'h01,8'h21,8'h26,8'h27,8'h27,8'h27,8'h24,8'h2c,8'h4e,8'h4f,8'hb3,8'hd1,8'hc4,8'h7c,8'h43,8'h62,8'h2f,8'h09,8'h26,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h23,8'h02,8'h00,8'h00,8'h3f,8'h6e,8'h79,8'h69,8'h59,8'h65,8'h82,8'h99,8'ha5,8'hab,8'hc2,8'hcc,8'hd0,8'hce,8'hcb,8'hcb,8'hcc,8'hc0,8'haa,8'h9b,8'h8d,8'h70,8'h57,8'h6b,8'h94,8'hb7,8'hcc,8'hcc,8'hc1,8'h84,8'h4c,8'h4b,8'h5e,8'h5f,8'h41,8'h14,8'h00,8'h00,8'h32,8'h26,8'h38,8'h24,8'h22,8'h26,8'h45,8'h2e,8'h2b,8'h24,8'h24,8'h29,8'h34,8'h2a,8'h23,8'h10,8'h00,8'h00,8'h00,8'h43,8'h55,8'h49,8'h43,8'h34,8'h43,8'h4b,8'h64,8'hb7,8'hc9,8'hca,8'hcb,8'hc9,8'hc8,8'hc8,8'ha8,8'h42,8'h56,8'h20,8'h00,8'h1a,8'h21,8'h24,8'h24,8'h23,8'h23,8'h24,8'h25,8'h22,8'h28,8'h42,8'h48,8'h37,8'h34,8'h35,8'h2f,8'h28,8'h31,8'h33,8'h33,8'h2d,8'h22,8'h24,8'h38,8'h39,8'h29,8'h23,8'h26,8'h23,8'h23,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h2b,8'h27,8'h21,8'h22,8'h60,8'hcd,8'hed,8'h86,8'h29,8'h2b,8'h40,8'h63,8'h9d,8'he5,8'hee,8'hac,8'h61,8'h48,8'h73,8'h53,8'h2c,8'h22,8'h22,8'h23,8'h25,8'h3c,8'h34,8'h2c,8'h39,8'h33,8'h26,8'h33,8'h3c,8'h45,8'h2f,8'h25,8'h11,8'h00,8'h20,8'h3a,8'h5c,8'h58,8'h63,8'h82,8'h8c,8'ha7,8'hc4,8'hc9,8'hc9,8'hc6,8'ha2,8'h60,8'h57,8'h5b,8'h2f,8'h00,8'h21,8'h26,8'h27,8'h27,8'h27,8'h27,8'h25,8'h22,8'h4c,8'h45,8'h85,8'hc8,8'hcc,8'h8b,8'h45,8'h60,8'h38,8'h16,8'h26,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h24,8'h1b,8'h00,8'h00,8'h2e,8'h6e,8'h8d,8'h71,8'h4d,8'h5a,8'h8e,8'hbb,8'hcb,8'hcf,8'hcc,8'hc4,8'hae,8'h92,8'h7e,8'h6b,8'h55,8'h51,8'h9f,8'hd3,8'hd1,8'hcf,8'hcc,8'hbe,8'ha5,8'hb8,8'hcb,8'hcc,8'hc6,8'hab,8'h68,8'h3b,8'h51,8'h6e,8'h51,8'h1c,8'h00,8'h00,8'h00,8'h24,8'h38,8'h28,8'h23,8'h22,8'h22,8'h2b,8'h5c,8'h32,8'h2a,8'h28,8'h2e,8'h2a,8'h22,8'h21,8'h00,8'h00,8'h00,8'h00,8'h19,8'h48,8'h4c,8'h49,8'h4d,8'h51,8'h55,8'h56,8'h34,8'h81,8'hca,8'hcb,8'hcc,8'hc9,8'hc9,8'hc7,8'hab,8'h44,8'h5c,8'h24,8'h00,8'h1c,8'h21,8'h23,8'h23,8'h23,8'h23,8'h23,8'h23,8'h24,8'h2c,8'h3b,8'h60,8'h30,8'h2b,8'h33,8'h3d,8'h34,8'h38,8'h45,8'h36,8'h36,8'h20,8'h1e,8'h26,8'h27,8'h23,8'h24,8'h24,8'h24,8'h24,8'h25,8'h25,8'h24,8'h23,8'h24,8'h26,8'h31,8'h27,8'h2c,8'h25,8'h20,8'h4b,8'hc8,8'hf8,8'had,8'h2f,8'h1e,8'h25,8'h26,8'h28,8'h5a,8'hd6,8'he5,8'h7d,8'h32,8'h2b,8'h3b,8'h2e,8'h24,8'h21,8'h23,8'h26,8'h27,8'h2d,8'h38,8'h29,8'h27,8'h30,8'h25,8'h27,8'h2e,8'h32,8'h2d,8'h37,8'h30,8'h29,8'h03,8'h00,8'h27,8'h4b,8'h49,8'h51,8'h8d,8'hc2,8'hc9,8'hc7,8'hc8,8'ha6,8'h51,8'h54,8'h5e,8'h22,8'h00,8'h20,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h20,8'h34,8'h4e,8'h5d,8'hbb,8'hce,8'ha0,8'h45,8'h62,8'h4a,8'h00,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h23,8'h00,8'h00,8'h28,8'h53,8'h7a,8'h82,8'h6c,8'h62,8'h95,8'hc2,8'hcc,8'hc0,8'ha4,8'h95,8'h7e,8'h68,8'h58,8'h46,8'h47,8'h51,8'h50,8'h30,8'h8d,8'hd6,8'hd0,8'hcf,8'hcc,8'hcc,8'hc9,8'hc8,8'hc7,8'hab,8'h83,8'h56,8'h4a,8'h62,8'h60,8'h33,8'h00,8'h00,8'h00,8'h18,8'h21,8'h26,8'h22,8'h24,8'h23,8'h24,8'h24,8'h28,8'h2d,8'h25,8'h3d,8'h40,8'h3d,8'h2c,8'h35,8'h23,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h33,8'h41,8'h65,8'hc7,8'hcf,8'hce,8'hcb,8'hc6,8'hc7,8'hac,8'h45,8'h62,8'h27,8'h00,8'h1e,8'h22,8'h24,8'h24,8'h24,8'h28,8'h28,8'h2a,8'h35,8'h41,8'h41,8'h40,8'h24,8'h2b,8'h35,8'h26,8'h2e,8'h35,8'h26,8'h26,8'h33,8'h23,8'h19,8'h20,8'h24,8'h25,8'h23,8'h23,8'h24,8'h26,8'h26,8'h26,8'h25,8'h24,8'h26,8'h29,8'h2a,8'h2e,8'h2a,8'h25,8'h55,8'hc5,8'hf5,8'hc2,8'h47,8'h22,8'h24,8'h24,8'h22,8'h22,8'h39,8'h78,8'h8f,8'h4e,8'h2b,8'h20,8'h20,8'h22,8'h25,8'h26,8'h2c,8'h42,8'h2d,8'h41,8'h49,8'h2c,8'h27,8'h29,8'h22,8'h26,8'h26,8'h2b,8'h30,8'h52,8'h46,8'h49,8'h3b,8'h17,8'h00,8'h00,8'h35,8'h46,8'h43,8'h6a,8'h9a,8'hb5,8'hbf,8'h5f,8'h36,8'h80,8'h52,8'h00,8'h23,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h25,8'h28,8'h4f,8'h51,8'h9e,8'hce,8'haa,8'h55,8'h4c,8'h52,8'h01,8'h23,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h24,8'h1b,8'h00,8'h00,8'h4b,8'h7e,8'h69,8'h62,8'h86,8'hb4,8'hc7,8'hd2,8'hbd,8'h88,8'h57,8'h45,8'h5c,8'h6b,8'h72,8'h7a,8'h6e,8'h5b,8'h67,8'h71,8'h55,8'hb0,8'hd2,8'hce,8'hca,8'hc8,8'hc5,8'hc7,8'hbe,8'h81,8'h43,8'h4c,8'h6c,8'h62,8'h31,8'h00,8'h00,8'h08,8'h1f,8'h22,8'h28,8'h24,8'h23,8'h22,8'h23,8'h22,8'h24,8'h26,8'h2b,8'h28,8'h26,8'h3c,8'h37,8'h42,8'h35,8'h3c,8'h34,8'h25,8'h18,8'h42,8'h38,8'h0b,8'h07,8'h1c,8'h20,8'h03,8'h00,8'h00,8'h04,8'h40,8'h69,8'hcf,8'hd3,8'hcc,8'hcb,8'hca,8'hcb,8'haa,8'h44,8'h63,8'h28,8'h00,8'h24,8'h28,8'h27,8'h2b,8'h3a,8'h39,8'h3f,8'h44,8'h49,8'h4a,8'h4c,8'h41,8'h24,8'h24,8'h24,8'h23,8'h25,8'h27,8'h23,8'h23,8'h24,8'h24,8'h17,8'h0d,8'h21,8'h26,8'h24,8'h24,8'h26,8'h26,8'h25,8'h27,8'h3c,8'h3e,8'h42,8'h40,8'h32,8'h2f,8'h24,8'h62,8'hd6,8'hf7,8'hcc,8'h4d,8'h22,8'h27,8'h25,8'h24,8'h24,8'h26,8'h23,8'h37,8'h58,8'h23,8'h24,8'h21,8'h22,8'h23,8'h28,8'h2c,8'h33,8'h51,8'h29,8'h26,8'h28,8'h23,8'h23,8'h23,8'h22,8'h27,8'h2e,8'h27,8'h26,8'h34,8'h2b,8'h26,8'h25,8'h23,8'h21,8'h20,8'h14,8'h00,8'h26,8'h43,8'h4c,8'h56,8'h87,8'h6b,8'h38,8'h59,8'h89,8'h63,8'h2f,8'h26,8'h27,8'h27,8'h27,8'h27,8'h26,8'h20,8'h49,8'h45,8'h83,8'hcc,8'hb3,8'h54,8'h50,8'h58,8'h07,8'h24,8'h28,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h23,8'h00,8'h00,8'h00,8'h60,8'h7c,8'h5a,8'h6b,8'ha6,8'hce,8'hd9,8'hc3,8'h8d,8'h54,8'h45,8'h57,8'h6e,8'h71,8'h5c,8'h42,8'h28,8'h00,8'h00,8'h27,8'h5a,8'h67,8'hc4,8'hcf,8'hc7,8'hc5,8'hc8,8'hca,8'hb0,8'h69,8'h36,8'h50,8'h6f,8'h47,8'h00,8'h00,8'h00,8'h16,8'h21,8'h26,8'h32,8'h38,8'h26,8'h22,8'h23,8'h25,8'h30,8'h2b,8'h2b,8'h28,8'h27,8'h29,8'h29,8'h25,8'h30,8'h2c,8'h52,8'h52,8'h55,8'h2e,8'h49,8'h43,8'h23,8'h2c,8'h32,8'h2f,8'h28,8'h19,8'h00,8'h05,8'h40,8'h71,8'hcf,8'hd0,8'hce,8'hce,8'hcd,8'hce,8'ha9,8'h43,8'h63,8'h25,8'h29,8'h5a,8'h38,8'h4f,8'h39,8'h3c,8'h54,8'h46,8'h33,8'h37,8'h3d,8'h4a,8'h34,8'h21,8'h23,8'h23,8'h24,8'h23,8'h23,8'h24,8'h25,8'h24,8'h23,8'h1e,8'h10,8'h20,8'h26,8'h2b,8'h2b,8'h26,8'h20,8'h21,8'h30,8'h53,8'h5f,8'h4a,8'h41,8'h28,8'h20,8'h53,8'hd0,8'hfb,8'he2,8'h67,8'h21,8'h23,8'h24,8'h24,8'h24,8'h24,8'h27,8'h27,8'h38,8'h57,8'h24,8'h27,8'h23,8'h26,8'h28,8'h29,8'h26,8'h25,8'h27,8'h22,8'h23,8'h24,8'h24,8'h24,8'h23,8'h23,8'h24,8'h26,8'h24,8'h24,8'h24,8'h24,8'h23,8'h24,8'h26,8'h23,8'h24,8'h25,8'h23,8'h00,8'h00,8'h35,8'h45,8'h45,8'h67,8'h78,8'h46,8'h4b,8'h89,8'h74,8'h2c,8'h23,8'h27,8'h27,8'h25,8'h16,8'h33,8'h4b,8'h5e,8'hc5,8'hca,8'h65,8'h44,8'h64,8'h25,8'h09,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h00,8'h22,8'h00,8'h00,8'h19,8'h6a,8'h6f,8'h58,8'h88,8'hc6,8'hd6,8'hd2,8'ha2,8'h5e,8'h45,8'h5a,8'h75,8'h62,8'h3e,8'h03,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2d,8'h56,8'h80,8'hca,8'hd0,8'hca,8'hcb,8'hc8,8'h9b,8'h4f,8'h37,8'h66,8'h6b,8'h2e,8'h00,8'h00,8'h0d,8'h22,8'h20,8'h23,8'h2c,8'h36,8'h2e,8'h24,8'h22,8'h23,8'h2a,8'h5c,8'h31,8'h26,8'h23,8'h25,8'h2a,8'h24,8'h46,8'h4c,8'h33,8'h43,8'h3c,8'h41,8'h2b,8'h2a,8'h26,8'h43,8'h4c,8'h2b,8'h32,8'h36,8'h25,8'h00,8'h0e,8'h43,8'h75,8'hd5,8'hd0,8'hd0,8'hd1,8'hd3,8'hd0,8'had,8'h45,8'h62,8'h22,8'h25,8'h52,8'h33,8'h46,8'h3f,8'h30,8'h44,8'h3c,8'h3e,8'h43,8'h28,8'h30,8'h28,8'h29,8'h32,8'h23,8'h23,8'h23,8'h24,8'h25,8'h25,8'h25,8'h24,8'h22,8'h23,8'h4a,8'h47,8'h66,8'h47,8'h26,8'h17,8'h1c,8'h2e,8'h30,8'h31,8'h27,8'h26,8'h21,8'h49,8'hc3,8'hf9,8'hf1,8'h8d,8'h26,8'h22,8'h25,8'h24,8'h24,8'h24,8'h23,8'h2b,8'h41,8'h3c,8'h51,8'h26,8'h28,8'h26,8'h26,8'h2f,8'h4f,8'h30,8'h23,8'h22,8'h22,8'h23,8'h25,8'h24,8'h25,8'h24,8'h25,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h23,8'h25,8'h27,8'h33,8'h34,8'h2e,8'h22,8'h03,8'h00,8'h1a,8'h43,8'h43,8'h53,8'h79,8'h5a,8'h42,8'h7a,8'h7c,8'h39,8'h23,8'h26,8'h21,8'h22,8'h53,8'h47,8'hab,8'hd8,8'h7f,8'h3c,8'h65,8'h35,8'h0d,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h25,8'h02,8'h00,8'h2e,8'h69,8'h61,8'h61,8'ha4,8'hd0,8'hd3,8'hbf,8'h7e,8'h46,8'h53,8'h77,8'h65,8'h39,8'h00,8'h00,8'h00,8'h00,8'h11,8'h12,8'h00,8'h00,8'h42,8'h55,8'h93,8'hcb,8'hcb,8'hce,8'hc2,8'h84,8'h41,8'h47,8'h6d,8'h58,8'h05,8'h00,8'h00,8'h23,8'h28,8'h30,8'h23,8'h24,8'h23,8'h21,8'h24,8'h24,8'h23,8'h25,8'h24,8'h2a,8'h2c,8'h24,8'h24,8'h24,8'h24,8'h2f,8'h54,8'h41,8'h32,8'h3f,8'h30,8'h2a,8'h28,8'h28,8'h27,8'h29,8'h41,8'h2b,8'h3d,8'h60,8'h2d,8'h00,8'h1f,8'h42,8'h75,8'hd5,8'hd1,8'hd3,8'hd4,8'hd3,8'hd0,8'hb1,8'h47,8'h60,8'h20,8'h29,8'h48,8'h2f,8'h2b,8'h40,8'h39,8'h35,8'h37,8'h65,8'h41,8'h23,8'h2d,8'h3c,8'h4b,8'h4e,8'h25,8'h24,8'h28,8'h26,8'h24,8'h24,8'h25,8'h26,8'h29,8'h26,8'h5f,8'h6a,8'h4a,8'h3e,8'h26,8'h15,8'h15,8'h25,8'h26,8'h24,8'h26,8'h24,8'h47,8'hc3,8'hf8,8'hf8,8'hba,8'h37,8'h21,8'h25,8'h25,8'h25,8'h25,8'h25,8'h24,8'h25,8'h33,8'h35,8'h42,8'h25,8'h24,8'h26,8'h24,8'h26,8'h2c,8'h26,8'h22,8'h23,8'h2a,8'h2b,8'h24,8'h23,8'h24,8'h25,8'h24,8'h25,8'h23,8'h24,8'h25,8'h25,8'h26,8'h25,8'h26,8'h2f,8'h2d,8'h3c,8'h50,8'h26,8'h21,8'h22,8'h20,8'h00,8'h00,8'h36,8'h48,8'h47,8'h6e,8'h63,8'h42,8'h68,8'h84,8'h49,8'h26,8'h20,8'h4b,8'h46,8'h7e,8'hd1,8'h9c,8'h42,8'h60,8'h51,8'h03,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h22,8'h00,8'h00,8'h2e,8'h6b,8'h5a,8'h6c,8'hbb,8'hd6,8'hd1,8'hae,8'h66,8'h47,8'h6a,8'h75,8'h47,8'h00,8'h00,8'h00,8'h06,8'h1c,8'h20,8'h23,8'h21,8'h00,8'h00,8'h4a,8'h5a,8'hac,8'hd0,8'hcc,8'hbb,8'h6e,8'h3f,8'h55,8'h6c,8'h44,8'h00,8'h00,8'h00,8'h2f,8'h42,8'h25,8'h2c,8'h23,8'h2c,8'h26,8'h21,8'h24,8'h26,8'h23,8'h28,8'h28,8'h21,8'h2b,8'h25,8'h22,8'h22,8'h22,8'h29,8'h3c,8'h2d,8'h27,8'h41,8'h36,8'h3f,8'h32,8'h27,8'h26,8'h2b,8'h53,8'h2e,8'h2f,8'h42,8'h26,8'h00,8'h1f,8'h3e,8'h76,8'hd4,8'hd3,8'hd3,8'hd6,8'hd3,8'hce,8'hac,8'h46,8'h61,8'h24,8'h23,8'h3c,8'h29,8'h27,8'h27,8'h28,8'h23,8'h25,8'h2d,8'h25,8'h28,8'h2a,8'h45,8'h49,8'h36,8'h21,8'h2e,8'h4a,8'h43,8'h23,8'h24,8'h25,8'h25,8'h30,8'h32,8'h43,8'h9a,8'h4d,8'h2b,8'h25,8'h27,8'h2f,8'h25,8'h26,8'h26,8'h26,8'h44,8'hb3,8'hf5,8'hf9,8'hd7,8'h55,8'h23,8'h27,8'h26,8'h26,8'h26,8'h26,8'h26,8'h29,8'h24,8'h2a,8'h36,8'h33,8'h24,8'h23,8'h23,8'h24,8'h23,8'h21,8'h26,8'h34,8'h22,8'h34,8'h3a,8'h23,8'h22,8'h23,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h26,8'h25,8'h29,8'h2c,8'h2a,8'h40,8'h49,8'h3c,8'h30,8'h3f,8'h2d,8'h3d,8'h2e,8'h0c,8'h00,8'h1c,8'h3d,8'h44,8'h5d,8'h69,8'h46,8'h58,8'h88,8'h61,8'h4e,8'h4d,8'h5c,8'hc2,8'haf,8'h4f,8'h58,8'h62,8'h18,8'h26,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h22,8'h00,8'h00,8'h45,8'h64,8'h6c,8'h88,8'hc7,8'hd1,8'hc4,8'h93,8'h5a,8'h52,8'h63,8'h51,8'h17,8'h00,8'h00,8'h0b,8'h1f,8'h21,8'h21,8'h22,8'h24,8'h21,8'h00,8'h00,8'h56,8'h6d,8'hc7,8'hc7,8'h9b,8'h62,8'h48,8'h5b,8'h58,8'h26,8'h00,8'h00,8'h13,8'h24,8'h42,8'h4a,8'h2e,8'h45,8'h2b,8'h24,8'h22,8'h26,8'h36,8'h2c,8'h23,8'h28,8'h34,8'h49,8'h28,8'h21,8'h28,8'h45,8'h42,8'h4e,8'h30,8'h26,8'h2a,8'h3f,8'h3e,8'h54,8'h30,8'h24,8'h24,8'h25,8'h29,8'h23,8'h22,8'h21,8'h17,8'h00,8'h21,8'h3f,8'h7e,8'hd6,8'hd4,8'hd1,8'hd5,8'hd1,8'hd0,8'had,8'h47,8'h62,8'h24,8'h20,8'h2c,8'h21,8'h22,8'h23,8'h24,8'h23,8'h27,8'h30,8'h26,8'h39,8'h45,8'h42,8'h2d,8'h2c,8'h2e,8'h3d,8'h43,8'h39,8'h22,8'h23,8'h24,8'h29,8'h36,8'h3a,8'h28,8'h82,8'hab,8'h44,8'h20,8'h36,8'h69,8'h2f,8'h21,8'h24,8'h4a,8'had,8'hf3,8'hf8,8'hd9,8'h6a,8'h24,8'h26,8'h28,8'h29,8'h2a,8'h29,8'h24,8'h26,8'h2b,8'h3a,8'h33,8'h2b,8'h26,8'h23,8'h23,8'h24,8'h22,8'h26,8'h2b,8'h32,8'h48,8'h24,8'h24,8'h28,8'h28,8'h24,8'h22,8'h22,8'h24,8'h24,8'h24,8'h2b,8'h4a,8'h2d,8'h24,8'h29,8'h42,8'h37,8'h3d,8'h49,8'h26,8'h2f,8'h41,8'h27,8'h43,8'h3f,8'h2e,8'h20,8'h0f,8'h07,8'h30,8'h3c,8'h53,8'h58,8'h4d,8'h53,8'h6c,8'h5a,8'h54,8'haa,8'hb1,8'h58,8'h4f,8'h5f,8'h23,8'h22,8'h2a,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h03,8'h00,8'h48,8'h66,8'h63,8'ha9,8'hd1,8'hd4,8'hc4,8'h84,8'h46,8'h65,8'h6b,8'h2b,8'h00,8'h00,8'h0e,8'h20,8'h21,8'h22,8'h21,8'h20,8'h28,8'h2b,8'h20,8'h00,8'h28,8'h55,8'h84,8'hc9,8'h80,8'h3e,8'h50,8'h6a,8'h3c,8'h00,8'h00,8'h07,8'h1f,8'h21,8'h24,8'h49,8'h4a,8'h2c,8'h4b,8'h2d,8'h16,8'h12,8'h2d,8'h57,8'h2e,8'h22,8'h26,8'h31,8'h57,8'h2e,8'h28,8'h33,8'h6f,8'hb8,8'hca,8'h68,8'h28,8'h27,8'h38,8'h2d,8'h25,8'h23,8'h22,8'h24,8'h24,8'h21,8'h22,8'h22,8'h24,8'h21,8'h00,8'h20,8'h40,8'h86,8'hd7,8'hd8,8'hd7,8'hd5,8'hd4,8'hd4,8'hb2,8'h4b,8'h67,8'h25,8'h03,8'h21,8'h22,8'h22,8'h23,8'h24,8'h24,8'h26,8'h29,8'h24,8'h30,8'h4b,8'h39,8'h35,8'h3e,8'h40,8'h28,8'h24,8'h24,8'h27,8'h27,8'h29,8'h2e,8'h40,8'h2e,8'h22,8'h43,8'hcc,8'ha4,8'h26,8'h2f,8'h95,8'h49,8'h1c,8'h4a,8'hc1,8'hf6,8'hfa,8'he8,8'h74,8'h23,8'h22,8'h29,8'h2f,8'h32,8'h2b,8'h31,8'h2e,8'h26,8'h24,8'h2e,8'h27,8'h22,8'h27,8'h36,8'h56,8'h30,8'h23,8'h29,8'h33,8'h29,8'h2a,8'h22,8'h22,8'h24,8'h25,8'h24,8'h22,8'h22,8'h21,8'h22,8'h23,8'h2b,8'h4b,8'h2f,8'h2b,8'h26,8'h34,8'h34,8'h24,8'h26,8'h2c,8'h21,8'h23,8'h2c,8'h33,8'h36,8'h52,8'h37,8'h51,8'h29,8'h00,8'h00,8'h37,8'h41,8'h48,8'h53,8'h35,8'h45,8'ha5,8'hc1,8'h56,8'h49,8'h61,8'h20,8'h22,8'h28,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h20,8'h00,8'h44,8'h65,8'h61,8'hb1,8'hd4,8'hce,8'hc8,8'h8b,8'h48,8'h64,8'h64,8'h25,8'h00,8'h00,8'h1e,8'h22,8'h23,8'h24,8'h25,8'h28,8'h32,8'h26,8'h24,8'h0b,8'h00,8'h43,8'h4c,8'h86,8'h79,8'h3a,8'h59,8'h64,8'h2b,8'h00,8'h00,8'h0f,8'h20,8'h21,8'h24,8'h27,8'h3b,8'h31,8'h21,8'h20,8'h07,8'h00,8'h22,8'h2b,8'h29,8'h29,8'h23,8'h26,8'h2b,8'h53,8'h2e,8'h28,8'h42,8'h7b,8'he2,8'hee,8'h91,8'h3b,8'h2a,8'h32,8'h27,8'h22,8'h23,8'h23,8'h21,8'h23,8'h24,8'h25,8'h26,8'h2a,8'h23,8'h00,8'h29,8'h45,8'h93,8'hd6,8'hd9,8'hda,8'hd5,8'hd6,8'hd1,8'hb3,8'h4d,8'h6c,8'h27,8'h02,8'h23,8'h21,8'h22,8'h29,8'h26,8'h24,8'h23,8'h24,8'h26,8'h2c,8'h29,8'h36,8'h37,8'h25,8'h24,8'h24,8'h23,8'h32,8'h55,8'h3e,8'h32,8'h46,8'h62,8'h2f,8'h23,8'h25,8'h96,8'he7,8'h6d,8'h37,8'hab,8'h6e,8'h43,8'hbd,8'hf7,8'hf9,8'hf0,8'h9b,8'h2c,8'h24,8'h2d,8'h2b,8'h29,8'h26,8'h25,8'h45,8'h46,8'h24,8'h23,8'h24,8'h25,8'h27,8'h2c,8'h39,8'h64,8'h31,8'h28,8'h26,8'h36,8'h35,8'h21,8'h21,8'h24,8'h21,8'h22,8'h21,8'h22,8'h1d,8'h11,8'h26,8'h26,8'h26,8'h25,8'h24,8'h26,8'h24,8'h24,8'h24,8'h23,8'h25,8'h2b,8'h24,8'h23,8'h39,8'h50,8'h28,8'h2b,8'h2a,8'h41,8'h2c,8'h23,8'h0a,8'h00,8'h2b,8'h41,8'h40,8'h69,8'h9e,8'hbe,8'h6f,8'h48,8'h68,8'h2d,8'h16,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h24,8'h09,8'h00,8'h4b,8'h61,8'h74,8'hb0,8'hd4,8'hd1,8'hc4,8'h81,8'h51,8'h6b,8'h64,8'h1c,8'h00,8'h0e,8'h21,8'h22,8'h23,8'h24,8'h25,8'h26,8'h45,8'h4c,8'h2e,8'h22,8'h00,8'h00,8'h54,8'h33,8'h4a,8'h52,8'h62,8'h4f,8'h20,8'h00,8'h35,8'h2c,8'h1a,8'h22,8'h24,8'h24,8'h24,8'h23,8'h1a,8'h00,8'h00,8'h00,8'h00,8'h30,8'h35,8'h23,8'h26,8'h24,8'h26,8'h26,8'h2d,8'h26,8'h22,8'h26,8'h48,8'h89,8'hac,8'h62,8'h28,8'h22,8'h23,8'h22,8'h22,8'h24,8'h23,8'h23,8'h22,8'h2c,8'h31,8'h36,8'h38,8'h23,8'h00,8'h2d,8'h45,8'h95,8'hd7,8'hd9,8'hd5,8'hd4,8'hcf,8'hd0,8'hb3,8'h4c,8'h69,8'h22,8'h1f,8'h3c,8'h2c,8'h2b,8'h2b,8'h28,8'h26,8'h2d,8'h2c,8'h28,8'h27,8'h25,8'h2f,8'h32,8'h23,8'h22,8'h24,8'h24,8'h39,8'h62,8'h40,8'h32,8'h35,8'h3e,8'h29,8'h25,8'h22,8'h4b,8'hd4,8'hd7,8'h96,8'hd1,8'hca,8'hbe,8'hf2,8'hf8,8'hf3,8'ha1,8'h36,8'h21,8'h22,8'h26,8'h26,8'h1e,8'h19,8'h25,8'h3a,8'h35,8'h23,8'h22,8'h25,8'h2b,8'h3f,8'h2e,8'h31,8'h33,8'h2e,8'h46,8'h24,8'h31,8'h2f,8'h22,8'h22,8'h21,8'h20,8'h1f,8'h0f,8'h00,8'h00,8'h00,8'h3b,8'h2b,8'h24,8'h24,8'h24,8'h25,8'h25,8'h24,8'h24,8'h25,8'h2e,8'h45,8'h27,8'h24,8'h28,8'h2f,8'h25,8'h26,8'h2b,8'h43,8'h45,8'h3f,8'h24,8'h00,8'h00,8'h4d,8'h3c,8'h8b,8'hc1,8'h68,8'h4e,8'h61,8'h32,8'h14,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h24,8'h00,8'h00,8'h46,8'h61,8'h68,8'hb6,8'hd8,8'hd8,8'hcd,8'h90,8'h46,8'h6f,8'h6e,8'h10,8'h00,8'h0c,8'h1f,8'h23,8'h23,8'h23,8'h24,8'h24,8'h24,8'h32,8'h3a,8'h51,8'h25,8'h00,8'h15,8'h4c,8'h1f,8'h46,8'h6c,8'h46,8'h00,8'h00,8'h12,8'h2f,8'h29,8'h21,8'h24,8'h29,8'h20,8'h06,8'h00,8'h00,8'h00,8'h00,8'h00,8'h16,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h23,8'h24,8'h24,8'h2c,8'h33,8'h37,8'h50,8'h34,8'h26,8'h23,8'h23,8'h23,8'h22,8'h24,8'h26,8'h24,8'h29,8'h52,8'h47,8'h46,8'h4a,8'h25,8'h00,8'h35,8'h49,8'h9b,8'hd9,8'hd9,8'hd7,8'hd9,8'hd3,8'hd1,8'hb3,8'h4c,8'h69,8'h1a,8'h12,8'h49,8'h48,8'h39,8'h24,8'h26,8'h28,8'h2c,8'h27,8'h28,8'h27,8'h25,8'h24,8'h23,8'h2c,8'h34,8'h31,8'h2c,8'h38,8'h68,8'h4e,8'h2e,8'h24,8'h23,8'h25,8'h24,8'h24,8'h22,8'h8c,8'hf5,8'hf4,8'hf5,8'hf8,8'hf9,8'hf7,8'hf8,8'hcb,8'h42,8'h23,8'h41,8'h5a,8'h51,8'h22,8'h0d,8'h1c,8'h26,8'h26,8'h24,8'h26,8'h26,8'h30,8'h2f,8'h3a,8'h2e,8'h2e,8'h2b,8'h28,8'h33,8'h27,8'h25,8'h23,8'h22,8'h1f,8'h13,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0d,8'h25,8'h24,8'h26,8'h24,8'h24,8'h25,8'h24,8'h25,8'h40,8'h39,8'h33,8'h56,8'h27,8'h24,8'h24,8'h27,8'h2b,8'h27,8'h27,8'h31,8'h3a,8'h31,8'h21,8'h00,8'h3a,8'h47,8'h5e,8'hb6,8'h6c,8'h46,8'h6c,8'h2d,8'h03,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h20,8'h00,8'h35,8'h66,8'h63,8'hb1,8'hd8,8'hd6,8'hd3,8'hae,8'h53,8'h66,8'h78,8'h2b,8'h00,8'h0a,8'h1f,8'h22,8'h24,8'h25,8'h23,8'h29,8'h2b,8'h25,8'h23,8'h26,8'h30,8'h23,8'h00,8'h37,8'h4b,8'h4e,8'h66,8'h33,8'h00,8'h00,8'h12,8'h22,8'h24,8'h22,8'h21,8'h22,8'h0d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h29,8'h48,8'h27,8'h24,8'h25,8'h25,8'h24,8'h24,8'h25,8'h25,8'h24,8'h26,8'h25,8'h2e,8'h43,8'h24,8'h22,8'h24,8'h24,8'h26,8'h2b,8'h26,8'h25,8'h27,8'h35,8'h3f,8'h2d,8'h40,8'h47,8'h21,8'h00,8'h37,8'h4a,8'ha8,8'hda,8'hd8,8'hd8,8'hd7,8'hd5,8'hd1,8'haf,8'h4b,8'h66,8'h0d,8'h00,8'h2a,8'h39,8'h2f,8'h30,8'h40,8'h26,8'h2c,8'h2f,8'h2d,8'h2f,8'h29,8'h26,8'h26,8'h48,8'h55,8'h30,8'h2b,8'h2e,8'h41,8'h37,8'h27,8'h28,8'h28,8'h28,8'h28,8'h28,8'h26,8'h62,8'he7,8'hf8,8'hf7,8'hf7,8'hf7,8'hf7,8'hf7,8'hd2,8'h91,8'h9c,8'ha8,8'h76,8'h3b,8'h21,8'h22,8'h24,8'h24,8'h26,8'h28,8'h2a,8'h2b,8'h26,8'h2b,8'h31,8'h2f,8'h24,8'h24,8'h26,8'h28,8'h3f,8'h22,8'h22,8'h13,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h21,8'h23,8'h25,8'h25,8'h26,8'h25,8'h26,8'h29,8'h42,8'h35,8'h2a,8'h3b,8'h28,8'h23,8'h2a,8'h29,8'h32,8'h2a,8'h26,8'h25,8'h25,8'h1f,8'h00,8'h1a,8'h4b,8'h49,8'h9a,8'h81,8'h45,8'h6e,8'h46,8'h00,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h23,8'h00,8'h40,8'h63,8'h66,8'hb7,8'hd5,8'hd0,8'hd0,8'hbb,8'h61,8'h65,8'h73,8'h2c,8'h00,8'h14,8'h22,8'h23,8'h24,8'h24,8'h24,8'h21,8'h35,8'h46,8'h4f,8'h2f,8'h27,8'h22,8'h06,8'h00,8'h55,8'h7e,8'h60,8'h1e,8'h00,8'h24,8'h25,8'h24,8'h22,8'h23,8'h1a,8'h00,8'h00,8'h00,8'h08,8'h47,8'h61,8'h47,8'h00,8'h00,8'h1a,8'h26,8'h2d,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h26,8'h26,8'h24,8'h22,8'h22,8'h30,8'h45,8'h23,8'h20,8'h22,8'h30,8'h5d,8'h4c,8'h43,8'h46,8'h48,8'h51,8'h42,8'h2a,8'h2c,8'h32,8'h20,8'h00,8'h3b,8'h4a,8'hab,8'hd8,8'hd5,8'hd9,8'hd8,8'hd5,8'hd2,8'hac,8'h48,8'h68,8'h23,8'h00,8'h21,8'h40,8'h50,8'h48,8'h44,8'h3a,8'h3e,8'h64,8'h41,8'h29,8'h2c,8'h25,8'h1c,8'h20,8'h24,8'h1b,8'h15,8'h27,8'h43,8'h56,8'h67,8'h80,8'h85,8'h87,8'h88,8'h8b,8'h9b,8'hbf,8'hf0,8'hf7,8'hf7,8'hf7,8'hf7,8'hf7,8'hf7,8'hf3,8'hb7,8'h61,8'h39,8'h24,8'h20,8'h23,8'h24,8'h27,8'h26,8'h35,8'h41,8'h4e,8'h4b,8'h22,8'h24,8'h28,8'h27,8'h22,8'h23,8'h21,8'h1f,8'h12,8'h00,8'h00,8'h00,8'h17,8'h48,8'h5a,8'h00,8'h00,8'h00,8'h1c,8'h22,8'h22,8'h24,8'h24,8'h26,8'h28,8'h27,8'h28,8'h2d,8'h2c,8'h24,8'h45,8'h57,8'h44,8'h25,8'h41,8'h31,8'h31,8'h2e,8'h27,8'h24,8'h26,8'h00,8'h13,8'h47,8'h4a,8'h8a,8'h6d,8'h47,8'h68,8'h40,8'h01,8'h24,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h21,8'h00,8'h24,8'h64,8'h60,8'ha7,8'hdd,8'hd9,8'hcd,8'hca,8'h7b,8'h4c,8'h83,8'h43,8'h00,8'h03,8'h22,8'h24,8'h23,8'h24,8'h25,8'h25,8'h22,8'h28,8'h3f,8'h4f,8'h45,8'h2a,8'h20,8'h00,8'h00,8'h6c,8'h67,8'h00,8'h00,8'h1f,8'h39,8'h25,8'h23,8'h0c,8'h00,8'h00,8'h00,8'h19,8'h43,8'h60,8'h82,8'h78,8'h16,8'h00,8'h0f,8'h23,8'h30,8'h32,8'h23,8'h24,8'h25,8'h24,8'h24,8'h24,8'h24,8'h25,8'h24,8'h1d,8'h0a,8'h01,8'h0f,8'h00,8'h00,8'h13,8'h28,8'h4f,8'h50,8'h5e,8'h52,8'h41,8'h35,8'h2f,8'h2b,8'h2e,8'h34,8'h21,8'h00,8'h3b,8'h46,8'hae,8'hd9,8'hd6,8'hd5,8'hd4,8'hd3,8'hd5,8'hab,8'h46,8'h6a,8'h24,8'h1f,8'h3f,8'h2e,8'h47,8'h4c,8'h46,8'h45,8'h40,8'h31,8'h28,8'h24,8'h25,8'h2d,8'h20,8'h1d,8'h1c,8'h19,8'h0d,8'h25,8'h42,8'h59,8'h75,8'h8f,8'hab,8'hc3,8'hd0,8'hdf,8'hed,8'hf7,8'hf7,8'hf7,8'hf7,8'hf7,8'hf7,8'hf8,8'hf9,8'hf6,8'ha0,8'h4b,8'h3b,8'h3d,8'h3c,8'h30,8'h24,8'h21,8'h22,8'h24,8'h22,8'h29,8'h2c,8'h22,8'h22,8'h22,8'h23,8'h17,8'h08,8'h00,8'h00,8'h00,8'h00,8'h26,8'h31,8'h40,8'h6d,8'h4e,8'h00,8'h00,8'h20,8'h22,8'h23,8'h22,8'h23,8'h24,8'h26,8'h2b,8'h2e,8'h4b,8'h3a,8'h2b,8'h24,8'h2d,8'h43,8'h41,8'h2c,8'h50,8'h4a,8'h30,8'h26,8'h23,8'h21,8'h08,8'h00,8'h4d,8'h41,8'h73,8'h72,8'h36,8'h62,8'h43,8'h00,8'h23,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h25,8'h00,8'h07,8'h60,8'h66,8'h96,8'hd8,8'hdc,8'hd8,8'hd2,8'ha2,8'h51,8'h72,8'h69,8'h00,8'h00,8'h20,8'h24,8'h25,8'h25,8'h24,8'h24,8'h23,8'h27,8'h3c,8'h43,8'h47,8'h35,8'h24,8'h20,8'h00,8'h00,8'h48,8'h06,8'h00,8'h20,8'h23,8'h1c,8'h13,8'h00,8'h00,8'h00,8'h24,8'h3a,8'h4f,8'h43,8'h3c,8'h6f,8'h4e,8'h00,8'h1a,8'h24,8'h28,8'h40,8'h40,8'h24,8'h22,8'h26,8'h26,8'h26,8'h21,8'h1a,8'h0d,8'h00,8'h00,8'h00,8'h00,8'h03,8'h01,8'h00,8'h00,8'h00,8'h00,8'h24,8'h2b,8'h2e,8'h28,8'h22,8'h24,8'h28,8'h4a,8'h4f,8'h25,8'h00,8'h3f,8'h47,8'hb1,8'hdb,8'hd8,8'hd8,8'hd7,8'hd5,8'hd7,8'hae,8'h47,8'h6c,8'h20,8'h16,8'h4c,8'h47,8'h42,8'h47,8'h4e,8'h42,8'h41,8'h28,8'h23,8'h24,8'h24,8'h29,8'h23,8'h21,8'h1b,8'h00,8'h00,8'h20,8'h2e,8'h3f,8'h44,8'h49,8'h51,8'h4b,8'h42,8'h5f,8'haf,8'hf2,8'hf8,8'hf7,8'hf7,8'hf7,8'hf7,8'hed,8'hd5,8'hc3,8'hac,8'h95,8'h89,8'h81,8'h76,8'h59,8'h2b,8'h17,8'h19,8'h19,8'h0e,8'h1c,8'h23,8'h21,8'h19,8'h09,8'h11,8'h00,8'h00,8'h11,8'h21,8'h35,8'h54,8'h56,8'h30,8'h41,8'h4c,8'h00,8'h00,8'h17,8'h22,8'h24,8'h33,8'h38,8'h31,8'h25,8'h26,8'h25,8'h25,8'h41,8'h44,8'h2e,8'h2e,8'h32,8'h28,8'h24,8'h2e,8'h2f,8'h46,8'h3d,8'h20,8'h19,8'h00,8'h00,8'h38,8'h47,8'h59,8'h72,8'h41,8'h6a,8'h77,8'h26,8'h00,8'h21,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h1b,8'h00,8'h5c,8'h66,8'h8a,8'hd8,8'hdf,8'hd8,8'hd6,8'hc5,8'h60,8'h63,8'h83,8'h24,8'h00,8'h1f,8'h24,8'h24,8'h25,8'h26,8'h25,8'h24,8'h26,8'h29,8'h28,8'h29,8'h2d,8'h24,8'h24,8'h1a,8'h00,8'h00,8'h00,8'h00,8'h04,8'h17,8'h00,8'h00,8'h00,8'h00,8'h35,8'h54,8'h47,8'h36,8'h40,8'h24,8'h4e,8'h5e,8'h00,8'h00,8'h43,8'h54,8'h3f,8'h37,8'h26,8'h24,8'h22,8'h25,8'h19,8'h00,8'h00,8'h00,8'h00,8'h15,8'h37,8'h56,8'h64,8'h68,8'h6a,8'h68,8'h5a,8'h31,8'h00,8'h00,8'h08,8'h20,8'h22,8'h23,8'h24,8'h28,8'h4e,8'h46,8'h21,8'h00,8'h3f,8'h45,8'hb6,8'hdc,8'hd5,8'hd9,8'hda,8'hd7,8'hdb,8'haf,8'h46,8'h68,8'h1c,8'h11,8'h41,8'h46,8'h39,8'h50,8'h5a,8'h4e,8'h2f,8'h27,8'h22,8'h22,8'h17,8'h00,8'h00,8'h00,8'h00,8'h2f,8'h53,8'h65,8'h5f,8'h5a,8'h56,8'h52,8'h41,8'h29,8'h44,8'h7a,8'hb1,8'he9,8'hf7,8'hf7,8'hf7,8'hf8,8'hf7,8'hae,8'h47,8'h33,8'h2e,8'h2c,8'h38,8'h49,8'h46,8'h3b,8'h2a,8'h24,8'h23,8'h22,8'h1a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1d,8'h3c,8'h4c,8'h49,8'h47,8'h69,8'h94,8'h6b,8'h4a,8'h4f,8'h00,8'h00,8'h00,8'h1e,8'h21,8'h24,8'h30,8'h50,8'h43,8'h22,8'h25,8'h27,8'h37,8'h39,8'h57,8'h32,8'h45,8'h44,8'h21,8'h22,8'h23,8'h21,8'h00,8'h00,8'h00,8'h00,8'h05,8'h40,8'h3f,8'h50,8'h62,8'h26,8'h30,8'h64,8'h85,8'h89,8'h58,8'h0e,8'h13,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h23,8'h00,8'h40,8'h6d,8'h71,8'hca,8'he0,8'hdb,8'hd8,8'hd6,8'ha0,8'h49,8'h81,8'h59,8'h00,8'h0b,8'h24,8'h26,8'h25,8'h26,8'h26,8'h26,8'h25,8'h29,8'h41,8'h2d,8'h24,8'h25,8'h22,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h14,8'h43,8'h54,8'h49,8'h3c,8'h4e,8'h84,8'h64,8'h33,8'h6e,8'h35,8'h00,8'h14,8'h28,8'h48,8'h33,8'h24,8'h21,8'h1d,8'h00,8'h00,8'h00,8'h00,8'h23,8'h3f,8'h50,8'h5b,8'h4f,8'h45,8'h3d,8'h3a,8'h3d,8'h42,8'h5b,8'h6c,8'h57,8'h12,8'h00,8'h06,8'h22,8'h24,8'h24,8'h25,8'h26,8'h25,8'h18,8'h00,8'h40,8'h46,8'hb9,8'hdc,8'hd7,8'hd9,8'hd7,8'hd8,8'hda,8'haf,8'h46,8'h67,8'h20,8'h23,8'h66,8'h43,8'h36,8'h40,8'h4e,8'h56,8'h24,8'h0a,8'h00,8'h00,8'h00,8'h00,8'h31,8'h4c,8'h5e,8'h67,8'h52,8'h45,8'h4b,8'h55,8'h50,8'h36,8'h2f,8'h35,8'h45,8'h3a,8'h46,8'hc0,8'hf9,8'hf9,8'hf7,8'hf9,8'hf8,8'h9e,8'h28,8'h22,8'h26,8'h2b,8'h32,8'h49,8'h55,8'h2b,8'h22,8'h19,8'h00,8'h00,8'h00,8'h00,8'h00,8'h19,8'h37,8'h49,8'h4e,8'h53,8'h5d,8'h7a,8'hac,8'hc7,8'h92,8'h4d,8'h5a,8'h20,8'h00,8'h00,8'h00,8'h04,8'h20,8'h23,8'h24,8'h28,8'h27,8'h24,8'h22,8'h2b,8'h50,8'h37,8'h2c,8'h28,8'h27,8'h27,8'h17,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2e,8'h4f,8'h64,8'h4f,8'h44,8'h80,8'h53,8'h4a,8'h59,8'h4e,8'h44,8'h5e,8'h90,8'h6e,8'h03,8'h09,8'h25,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h00,8'h27,8'h69,8'h6c,8'hb7,8'he2,8'hde,8'hd9,8'hd7,8'hcd,8'h6d,8'h63,8'h76,8'h22,8'h00,8'h1e,8'h24,8'h25,8'h26,8'h26,8'h26,8'h26,8'h26,8'h25,8'h2b,8'h28,8'h23,8'h24,8'h24,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2e,8'h3b,8'h41,8'h56,8'h61,8'h6d,8'h91,8'hc2,8'h9d,8'h40,8'h56,8'h52,8'h00,8'h00,8'h26,8'h20,8'h20,8'h19,8'h00,8'h00,8'h00,8'h07,8'h36,8'h39,8'h3a,8'h4c,8'h5e,8'h64,8'h71,8'h70,8'h72,8'h8b,8'h99,8'h99,8'h83,8'h6e,8'h59,8'h59,8'h64,8'h2b,8'h00,8'h11,8'h24,8'h26,8'h25,8'h24,8'h25,8'h17,8'h00,8'h40,8'h45,8'hb9,8'hde,8'hd9,8'hda,8'hd9,8'hd7,8'hd8,8'hb0,8'h48,8'h68,8'h0f,8'h11,8'h30,8'h29,8'h24,8'h18,8'h12,8'h00,8'h00,8'h05,8'h32,8'h44,8'h45,8'h46,8'h52,8'h63,8'h66,8'h6e,8'h71,8'h92,8'hbd,8'hce,8'hc8,8'hb0,8'hab,8'ha9,8'h8f,8'h40,8'h63,8'he1,8'he9,8'hba,8'hcf,8'hbe,8'he3,8'hb5,8'h35,8'h32,8'h3f,8'h34,8'h2b,8'h30,8'h24,8'h00,8'h00,8'h00,8'h00,8'h27,8'h32,8'h2d,8'h3a,8'h59,8'h6e,8'h7b,8'h7c,8'h9b,8'hc0,8'hd4,8'hd2,8'h9b,8'h51,8'h6b,8'h71,8'h45,8'h48,8'h50,8'h04,8'h00,8'h21,8'h23,8'h22,8'h23,8'h32,8'h47,8'h2b,8'h3f,8'h2f,8'h28,8'h24,8'h17,8'h03,8'h00,8'h00,8'h00,8'h23,8'h3f,8'h43,8'h46,8'h55,8'h64,8'h69,8'h72,8'h99,8'hbf,8'hb4,8'hc6,8'hc9,8'hc0,8'h99,8'h62,8'h57,8'h81,8'h65,8'h1c,8'h20,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h15,8'h00,8'h61,8'h5f,8'h96,8'hdb,8'hdd,8'hdb,8'hdb,8'hd5,8'hac,8'h4d,8'h82,8'h4f,8'h00,8'h12,8'h23,8'h26,8'h26,8'h26,8'h26,8'h27,8'h2b,8'h28,8'h23,8'h24,8'h24,8'h24,8'h26,8'h23,8'h07,8'h00,8'h00,8'h00,8'h00,8'h30,8'h4e,8'h46,8'h38,8'h51,8'h90,8'hbd,8'hcf,8'hd3,8'hc4,8'h5c,8'h46,8'h68,8'h0a,8'h00,8'h00,8'h03,8'h00,8'h00,8'h00,8'h00,8'h31,8'h4b,8'h4e,8'h47,8'h43,8'h56,8'h78,8'h9c,8'hba,8'hcd,8'hd4,8'hd4,8'hd7,8'hd7,8'hd6,8'hd4,8'hd0,8'ha3,8'h45,8'h52,8'h71,8'h0d,8'h00,8'h20,8'h24,8'h24,8'h26,8'h28,8'h0c,8'h00,8'h41,8'h50,8'hc2,8'hdb,8'hda,8'hdc,8'hdc,8'hd9,8'hda,8'hb0,8'h47,8'h65,8'h07,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2d,8'h50,8'h62,8'h5a,8'h47,8'h42,8'h4a,8'h6b,8'h97,8'hb6,8'hcc,8'hd1,8'hd5,8'hd6,8'hd7,8'hd9,8'hdc,8'hdc,8'hdc,8'ha5,8'h69,8'hd0,8'he6,8'h7b,8'h3a,8'h88,8'h60,8'ha5,8'hc1,8'h4c,8'h55,8'h35,8'h26,8'h06,8'h00,8'h00,8'h00,8'h29,8'h48,8'h4f,8'h45,8'h45,8'h59,8'h75,8'h9f,8'hba,8'hcc,8'hd2,8'hd5,8'hd7,8'hd8,8'hcc,8'h61,8'h33,8'h4f,8'h47,8'h43,8'h37,8'h64,8'h44,8'h00,8'h20,8'h22,8'h23,8'h24,8'h30,8'h44,8'h28,8'h35,8'h22,8'h00,8'h00,8'h00,8'h00,8'h17,8'h42,8'h5c,8'h61,8'h4d,8'h45,8'h53,8'h77,8'h9f,8'hc0,8'hd4,8'hd8,8'hd5,8'hd7,8'hd8,8'hd2,8'hd1,8'hd4,8'hc5,8'h6a,8'h44,8'h90,8'h4d,8'h01,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h22,8'h00,8'h45,8'h6d,8'h6a,8'hc9,8'hdb,8'hda,8'hd4,8'hd7,8'hd7,8'h83,8'h5a,8'h81,8'h28,8'h00,8'h21,8'h24,8'h25,8'h26,8'h26,8'h26,8'h27,8'h4f,8'h3c,8'h23,8'h25,8'h25,8'h23,8'h22,8'h03,8'h00,8'h00,8'h00,8'h21,8'h62,8'h53,8'h33,8'h4d,8'h86,8'hbc,8'hd6,8'hd4,8'hcf,8'hcc,8'h8e,8'h3b,8'h67,8'h42,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h44,8'h5a,8'h52,8'h42,8'h49,8'h6c,8'h9a,8'hbc,8'hce,8'hd7,8'hd4,8'hce,8'hce,8'hd3,8'hd3,8'hd5,8'hd1,8'hd1,8'hd4,8'hce,8'h8f,8'h3c,8'h6b,8'h50,8'h00,8'h11,8'h22,8'h23,8'h2d,8'h31,8'h0c,8'h00,8'h43,8'h53,8'hc4,8'hda,8'hd9,8'hdd,8'hdd,8'hdc,8'hdb,8'hb1,8'h4b,8'h6e,8'h22,8'h00,8'h00,8'h01,8'h35,8'h4d,8'h61,8'h61,8'h4f,8'h40,8'h48,8'h68,8'h90,8'hb4,8'hcc,8'hd4,8'hd4,8'hd5,8'hd3,8'hd2,8'hd5,8'hd5,8'hd3,8'hd6,8'hd5,8'hc5,8'h74,8'h9f,8'hd7,8'h7b,8'h3e,8'h22,8'h6b,8'h42,8'h5a,8'hbe,8'h55,8'h2f,8'h26,8'h01,8'h00,8'h11,8'h38,8'h56,8'h58,8'h48,8'h49,8'h68,8'h98,8'hbd,8'hca,8'hd2,8'hd2,8'hd2,8'hd3,8'hd0,8'hcf,8'hd4,8'hd3,8'h8a,8'h4c,8'h5d,8'h79,8'h8f,8'h54,8'h48,8'h44,8'h00,8'h1e,8'h22,8'h25,8'h22,8'h23,8'h21,8'h00,8'h00,8'h00,8'h00,8'h01,8'h34,8'h55,8'h6a,8'h64,8'h4c,8'h4a,8'h69,8'h96,8'hb5,8'hcd,8'hce,8'hce,8'hd3,8'hce,8'hcb,8'hcc,8'hd1,8'hd1,8'hd2,8'hd3,8'hd3,8'hae,8'h40,8'h73,8'h7b,8'h00,8'h24,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h25,8'h00,8'h26,8'h69,8'h66,8'hb1,8'hd8,8'hdb,8'hda,8'hd9,8'hd5,8'hb8,8'h55,8'h73,8'h67,8'h00,8'h0c,8'h24,8'h26,8'h27,8'h26,8'h33,8'h52,8'h2a,8'h38,8'h2c,8'h24,8'h27,8'h2b,8'h29,8'h38,8'h2f,8'h22,8'h00,8'h00,8'h13,8'h66,8'h5a,8'h40,8'ha6,8'hcd,8'hd0,8'hd5,8'hd2,8'hce,8'had,8'h4c,8'h52,8'h55,8'h00,8'h00,8'h2a,8'h3b,8'h33,8'h2e,8'h30,8'h46,8'h63,8'h83,8'h8e,8'hae,8'hcb,8'hd3,8'hd4,8'hd4,8'hd2,8'hcf,8'hce,8'hcd,8'hcd,8'hca,8'hcf,8'hcf,8'hcf,8'hd3,8'hd0,8'hca,8'h73,8'h50,8'h66,8'h00,8'h11,8'h30,8'h2b,8'h49,8'h37,8'h0b,8'h00,8'h47,8'h5d,8'hca,8'hda,8'hd9,8'hd9,8'hda,8'hd7,8'hd9,8'hae,8'h45,8'h83,8'h6b,8'h64,8'h5e,8'h4d,8'h43,8'h3c,8'h31,8'h47,8'h6b,8'h7f,8'ha4,8'hc4,8'hd4,8'hd6,8'hd4,8'hd4,8'hd4,8'hd3,8'hd2,8'hd4,8'hd0,8'hd0,8'hd1,8'hcf,8'hc8,8'h86,8'h88,8'ha1,8'h5a,8'h4c,8'h95,8'h35,8'h42,8'h37,8'h26,8'h7b,8'h55,8'h21,8'h16,8'h00,8'h43,8'h61,8'h4b,8'h66,8'h84,8'h97,8'hb3,8'hc9,8'hce,8'hcd,8'hcc,8'hcd,8'hcf,8'hcd,8'hcd,8'hcd,8'hd1,8'hd4,8'hd4,8'hc8,8'hbf,8'hc6,8'hd0,8'hcf,8'h70,8'h46,8'h44,8'h00,8'h1c,8'h1f,8'h05,8'h00,8'h00,8'h00,8'h00,8'h31,8'h4c,8'h52,8'h4d,8'h42,8'h48,8'h61,8'h80,8'h91,8'haf,8'hcc,8'hd2,8'hcf,8'hd2,8'hce,8'hca,8'hca,8'hcc,8'hcb,8'hcf,8'hce,8'hce,8'hcc,8'hcf,8'hd0,8'hcb,8'h67,8'h53,8'h94,8'h29,8'h21,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h1a,8'h00,8'h57,8'h60,8'h84,8'hda,8'hdb,8'hd7,8'hd9,8'hd7,8'hd4,8'h94,8'h4c,8'h86,8'h45,8'h00,8'h1b,8'h25,8'h26,8'h2f,8'h39,8'h35,8'h5c,8'h4b,8'h2a,8'h23,8'h27,8'h2b,8'h28,8'h2c,8'h37,8'h41,8'h42,8'h23,8'h00,8'h00,8'h00,8'h64,8'h4e,8'h83,8'hcd,8'hce,8'hd1,8'hce,8'hcb,8'h6e,8'h36,8'h7a,8'h60,8'h48,8'h67,8'h66,8'h45,8'h2d,8'h27,8'h24,8'h37,8'h56,8'h65,8'h66,8'h68,8'h7f,8'hc0,8'hd5,8'hd4,8'hd1,8'hcd,8'hd3,8'hce,8'hcc,8'hcb,8'hce,8'hd0,8'hce,8'hd0,8'hd0,8'hd5,8'h95,8'h45,8'h69,8'h00,8'h1c,8'h51,8'h41,8'h52,8'h3f,8'h00,8'h00,8'h48,8'h64,8'hcc,8'hd9,8'hda,8'hd7,8'hd7,8'hd6,8'hd8,8'ha8,8'h43,8'h8e,8'h9f,8'h93,8'h6b,8'h49,8'h38,8'h2f,8'h2e,8'h3b,8'h44,8'h4c,8'h52,8'h56,8'h80,8'hc7,8'hd6,8'hd4,8'hd6,8'hd4,8'hd0,8'hd3,8'hd0,8'hd4,8'hd3,8'hd0,8'h99,8'h65,8'h7d,8'h67,8'h5b,8'h5c,8'ha4,8'h35,8'h27,8'h27,8'h20,8'h46,8'h48,8'h20,8'h00,8'h0c,8'h61,8'h41,8'h6e,8'hb5,8'hd0,8'hd6,8'hd4,8'hcf,8'hcb,8'hca,8'hce,8'hce,8'hce,8'hce,8'hcd,8'hce,8'hce,8'hd0,8'hd1,8'hcd,8'hcd,8'hce,8'hce,8'hcd,8'h69,8'h4d,8'h3d,8'h00,8'h20,8'h14,8'h00,8'h00,8'h00,8'h00,8'h3e,8'h6e,8'h77,8'h50,8'h36,8'h27,8'h30,8'h4f,8'h61,8'h6c,8'h7c,8'h9c,8'hc8,8'hce,8'hcf,8'hce,8'hcf,8'hcb,8'hc9,8'hcc,8'hcb,8'hc9,8'hcd,8'hcd,8'hce,8'hcf,8'hd1,8'h82,8'h42,8'h90,8'h39,8'h21,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h24,8'h00,8'h2f,8'h6e,8'h61,8'hbc,8'hdd,8'hdb,8'hda,8'hd8,8'hd6,8'hce,8'h77,8'h58,8'h7e,8'h21,8'h00,8'h21,8'h27,8'h26,8'h36,8'h49,8'h2a,8'h2b,8'h3c,8'h27,8'h35,8'h40,8'h28,8'h2a,8'h3d,8'h46,8'h3c,8'h38,8'h2b,8'h23,8'h03,8'h00,8'h26,8'h58,8'h5e,8'hbf,8'hd6,8'hd2,8'hd4,8'hb4,8'h42,8'h59,8'h84,8'h6b,8'h63,8'h65,8'h59,8'h4d,8'h4f,8'h4d,8'h4d,8'h4b,8'h4c,8'h4c,8'h4b,8'h4d,8'h41,8'h73,8'hcf,8'hd4,8'hd3,8'hd0,8'hd0,8'hd0,8'hd1,8'hd3,8'hd5,8'hd1,8'hcf,8'hd0,8'hce,8'hd2,8'h96,8'h43,8'h67,8'h00,8'h20,8'h34,8'h2e,8'h45,8'h40,8'h00,8'h00,8'h48,8'h66,8'hcf,8'hda,8'hdb,8'hd9,8'hd4,8'hd7,8'hdb,8'haa,8'h43,8'h7c,8'h57,8'h44,8'h50,8'h54,8'h55,8'h59,8'h5c,8'h5b,8'h54,8'h51,8'h4a,8'h37,8'h30,8'h82,8'hd2,8'hd6,8'hd3,8'hd2,8'hd0,8'hd5,8'hd4,8'hd3,8'hd1,8'hb4,8'h4f,8'h47,8'h6e,8'hab,8'h80,8'h5e,8'h81,8'h01,8'h09,8'h1c,8'h23,8'h28,8'h27,8'h0c,8'h00,8'h3a,8'h53,8'h55,8'hbd,8'hd3,8'hd0,8'hd5,8'hd3,8'hd0,8'hd1,8'hce,8'hcf,8'hcf,8'hc7,8'hb8,8'ha5,8'h7e,8'h8d,8'hce,8'hd6,8'hd3,8'hd2,8'hd0,8'hce,8'hc6,8'h62,8'h57,8'h30,8'h00,8'h23,8'h19,8'h00,8'h00,8'h00,8'h00,8'h00,8'h11,8'h24,8'h29,8'h2f,8'h35,8'h3d,8'h41,8'h3f,8'h3c,8'h30,8'h42,8'h87,8'hca,8'hd2,8'hcf,8'hcc,8'hcb,8'hc8,8'hca,8'hc8,8'hcf,8'hcf,8'hcd,8'hd0,8'hd0,8'hcf,8'h8f,8'h41,8'h8b,8'h36,8'h20,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h1a,8'h06,8'h70,8'h55,8'h86,8'hdd,8'hda,8'hd8,8'hd5,8'hd5,8'hd6,8'hbd,8'h5c,8'h6f,8'h67,8'h00,8'h07,8'h3e,8'h39,8'h25,8'h2b,8'h2c,8'h29,8'h32,8'h2c,8'h28,8'h35,8'h32,8'h26,8'h2c,8'h2b,8'h3c,8'h42,8'h57,8'h2c,8'h24,8'h21,8'h00,8'h00,8'h4c,8'h53,8'h9b,8'hd9,8'hd6,8'hd3,8'hbd,8'h4c,8'h62,8'h69,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h42,8'h60,8'h46,8'hbc,8'hd5,8'hd3,8'hd4,8'hd2,8'hd2,8'hd1,8'hd0,8'hd5,8'hd4,8'hd0,8'hcf,8'hcd,8'hd1,8'h8e,8'h42,8'h66,8'h00,8'h21,8'h2a,8'h24,8'h3d,8'h37,8'h00,8'h00,8'h42,8'h62,8'hcf,8'hd9,8'hd9,8'hd9,8'hd7,8'hda,8'hdc,8'hab,8'h44,8'h6e,8'h15,8'h00,8'h10,8'h09,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h37,8'h4c,8'h48,8'hc0,8'hd8,8'hd6,8'hd6,8'hd8,8'hd6,8'hd4,8'hd7,8'hc6,8'h5e,8'h3c,8'h88,8'hc4,8'hd5,8'h70,8'h61,8'h5d,8'h00,8'h15,8'h44,8'h42,8'h22,8'h10,8'h00,8'h00,8'h54,8'h4a,8'h8f,8'hd6,8'hd7,8'hd6,8'hd7,8'hd5,8'hd4,8'hd6,8'hcf,8'hc1,8'h97,8'h60,8'h46,8'h40,8'h2b,8'h86,8'hd9,8'hd7,8'hd3,8'hd0,8'hd0,8'hcf,8'hbb,8'h50,8'h5f,8'h26,8'h00,8'h21,8'h25,8'h24,8'h25,8'h27,8'h2c,8'h1a,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h66,8'h4c,8'haf,8'hd1,8'hcd,8'hcb,8'hc8,8'hc8,8'hcc,8'hce,8'hcf,8'hcc,8'hce,8'hcd,8'hcd,8'hd2,8'h90,8'h3e,8'h8a,8'h35,8'h20,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h24,8'h00,8'h48,8'h75,8'h4a,8'hbb,8'he1,8'hda,8'hda,8'hd6,8'hd2,8'hd1,8'ha7,8'h49,8'h7c,8'h4c,8'h00,8'h1f,8'h46,8'h4e,8'h40,8'h31,8'h33,8'h32,8'h30,8'h2c,8'h2c,8'h2e,8'h26,8'h24,8'h27,8'h2a,8'h24,8'h2a,8'h30,8'h23,8'h24,8'h27,8'h1f,8'h00,8'h39,8'h4b,8'h81,8'hd1,8'hd7,8'hd5,8'hd0,8'h7a,8'h46,8'h72,8'h0e,8'h00,8'h00,8'h24,8'h29,8'h26,8'h11,8'h00,8'h00,8'h00,8'h00,8'h27,8'h5a,8'h4a,8'h5c,8'hc6,8'hd7,8'hd4,8'hd3,8'hcf,8'hce,8'hd0,8'hce,8'hd3,8'hd1,8'hd0,8'hd5,8'hd3,8'hd1,8'h8a,8'h41,8'h69,8'h05,8'h22,8'h2c,8'h2b,8'h46,8'h31,8'h00,8'h00,8'h3e,8'h61,8'hd0,8'hd8,8'hd8,8'hd9,8'hd8,8'hd8,8'hda,8'ha9,8'h46,8'h6d,8'h20,8'h21,8'h26,8'h26,8'h24,8'h21,8'h10,8'h00,8'h00,8'h00,8'h21,8'h53,8'h4b,8'h50,8'hc6,8'hd9,8'hd5,8'hd6,8'hd7,8'hd5,8'hd6,8'hd8,8'hac,8'h61,8'h9e,8'hd6,8'hda,8'hcf,8'h67,8'h65,8'h4f,8'h00,8'h0f,8'h2d,8'h38,8'h25,8'h25,8'h00,8'h00,8'h5e,8'h52,8'haf,8'hd9,8'hd4,8'hd7,8'hd7,8'hd7,8'hd6,8'hc3,8'h91,8'h5b,8'h3f,8'h44,8'h5c,8'h63,8'h38,8'haa,8'hdc,8'hd6,8'hd2,8'hd1,8'hd4,8'hd0,8'ha8,8'h4a,8'h65,8'h16,8'h02,8'h22,8'h49,8'h39,8'h34,8'h28,8'h2a,8'h24,8'h21,8'h25,8'h24,8'h25,8'h16,8'h00,8'h00,8'h00,8'h00,8'h4e,8'h7b,8'h4a,8'hb2,8'hd6,8'hce,8'hce,8'hc9,8'hcd,8'hd0,8'hd2,8'hcf,8'hcb,8'hcc,8'hcd,8'hcd,8'hd2,8'h8f,8'h40,8'h8c,8'h36,8'h20,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h0e,8'h00,8'h74,8'h51,8'h6d,8'hd4,8'hd9,8'hd5,8'hd6,8'hd5,8'hd1,8'hd0,8'h8c,8'h45,8'h7e,8'h36,8'h00,8'h22,8'h27,8'h41,8'h50,8'h57,8'h41,8'h2b,8'h28,8'h33,8'h2d,8'h2b,8'h27,8'h24,8'h25,8'h29,8'h26,8'h24,8'h23,8'h24,8'h2f,8'h30,8'h24,8'h00,8'h2e,8'h46,8'h7a,8'hd1,8'hd1,8'hd2,8'hd2,8'had,8'h46,8'h6f,8'h4c,8'h00,8'h14,8'h3a,8'h3b,8'h26,8'h00,8'h00,8'h00,8'h28,8'h49,8'h52,8'h45,8'h5a,8'haa,8'hd1,8'hd4,8'hd4,8'hd2,8'hce,8'hcd,8'hd3,8'hd4,8'hd4,8'hd2,8'hd5,8'hd4,8'hd1,8'hd0,8'h87,8'h44,8'h66,8'h00,8'h1e,8'h37,8'h3c,8'h2f,8'h26,8'h00,8'h00,8'h40,8'h64,8'hd5,8'hdb,8'hda,8'hdb,8'hd9,8'hdb,8'hdc,8'haa,8'h45,8'h70,8'h21,8'h23,8'h27,8'h27,8'h27,8'h27,8'h25,8'h00,8'h1f,8'h46,8'h53,8'h45,8'h41,8'h94,8'hd5,8'hd7,8'hd4,8'hd3,8'hd6,8'hd6,8'hd0,8'hd6,8'hcc,8'hc1,8'hd8,8'hdb,8'hda,8'hcf,8'h65,8'h69,8'h48,8'h00,8'h17,8'h21,8'h23,8'h23,8'h2f,8'h00,8'h23,8'h60,8'h59,8'hc2,8'hd9,8'hd6,8'hd6,8'hd5,8'hcf,8'ha3,8'h60,8'h44,8'h4a,8'h4e,8'h43,8'h3b,8'h5b,8'h41,8'hb7,8'hdc,8'hd7,8'hd5,8'hd3,8'hd4,8'hd2,8'h90,8'h48,8'h61,8'h00,8'h17,8'h23,8'h3a,8'h2f,8'h24,8'h23,8'h23,8'h23,8'h33,8'h4b,8'h37,8'h2d,8'h20,8'h00,8'h00,8'h31,8'h65,8'h6d,8'h44,8'h5d,8'hc6,8'hd4,8'hcd,8'hd2,8'hcb,8'hce,8'hca,8'hc6,8'hcd,8'hcd,8'hce,8'hd0,8'hd0,8'hd0,8'h88,8'h3f,8'h87,8'h31,8'h1f,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h23,8'h00,8'h3e,8'h77,8'h41,8'ha2,8'hde,8'hd7,8'hd7,8'hd7,8'hd7,8'hd5,8'hce,8'h75,8'h50,8'h7c,8'h1f,8'h00,8'h22,8'h25,8'h26,8'h36,8'h57,8'h3a,8'h24,8'h2f,8'h5b,8'h31,8'h23,8'h25,8'h24,8'h24,8'h24,8'h26,8'h2b,8'h3c,8'h46,8'h58,8'h33,8'h03,8'h00,8'h3f,8'h4a,8'h84,8'hd3,8'hd2,8'hd2,8'hd1,8'hcb,8'h66,8'h5b,8'h77,8'h00,8'h03,8'h48,8'h35,8'h22,8'h00,8'h00,8'h56,8'h62,8'h48,8'h54,8'h89,8'hc0,8'hd3,8'hd2,8'hce,8'hd0,8'hcd,8'hcd,8'hca,8'hb3,8'hae,8'hd2,8'hd4,8'hd5,8'hd2,8'hd2,8'hd5,8'h83,8'h46,8'h65,8'h00,8'h39,8'h57,8'h41,8'h42,8'h2c,8'h00,8'h00,8'h3d,8'h65,8'hd5,8'hdd,8'hdc,8'hdc,8'hdb,8'hdd,8'he0,8'had,8'h46,8'h6e,8'h1e,8'h23,8'h27,8'h27,8'h27,8'h25,8'h00,8'h3b,8'h5c,8'h4a,8'h3c,8'h5f,8'ha3,8'hd1,8'hd9,8'hd7,8'hd5,8'hd7,8'hc7,8'h96,8'h71,8'hbf,8'hdf,8'hdc,8'hdb,8'hdc,8'hde,8'hcc,8'h62,8'h6c,8'h43,8'h00,8'h21,8'h24,8'h22,8'h23,8'h22,8'h00,8'h3c,8'h57,8'h6d,8'hd5,8'hdb,8'hd9,8'hd8,8'hcd,8'h82,8'h45,8'h48,8'h51,8'h3d,8'h00,8'h00,8'h20,8'h4d,8'h4c,8'hc5,8'hde,8'hdc,8'hd6,8'hd6,8'hda,8'hd2,8'h72,8'h4c,8'h4f,8'h00,8'h21,8'h22,8'h22,8'h23,8'h24,8'h24,8'h23,8'h28,8'h37,8'h5c,8'h38,8'h1e,8'h00,8'h00,8'h53,8'h75,8'h56,8'h37,8'h58,8'hab,8'hcf,8'hca,8'hc7,8'hcb,8'hca,8'hbb,8'h81,8'h65,8'hb3,8'hca,8'hca,8'hcb,8'hce,8'hcc,8'h81,8'h41,8'h87,8'h2d,8'h1f,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h26,8'h14,8'h00,8'h68,8'h5a,8'h57,8'hcc,8'he0,8'hd8,8'hda,8'hdc,8'hdb,8'hd8,8'hd3,8'h69,8'h62,8'h7a,8'h00,8'h00,8'h29,8'h40,8'h3a,8'h2f,8'h45,8'h28,8'h24,8'h29,8'h38,8'h26,8'h23,8'h24,8'h24,8'h23,8'h24,8'h28,8'h34,8'h4f,8'h44,8'h50,8'h30,8'h00,8'h00,8'h50,8'h4d,8'ha0,8'hd7,8'hd7,8'hd6,8'hd4,8'hd4,8'h97,8'h48,8'h82,8'h43,8'h00,8'h2e,8'h37,8'h21,8'h00,8'h35,8'h64,8'h44,8'h81,8'hb7,8'hd0,8'hd5,8'hd1,8'hd2,8'hcc,8'hcd,8'hc9,8'hb3,8'h78,8'h3c,8'h65,8'hcb,8'hd0,8'hcf,8'hce,8'hd1,8'hd2,8'h7b,8'h4b,8'h62,8'h00,8'h37,8'h63,8'h46,8'h56,8'h30,8'h00,8'h00,8'h3f,8'h61,8'hc5,8'hce,8'hce,8'hcf,8'hce,8'hd0,8'hce,8'h9b,8'h46,8'h6c,8'h17,8'h24,8'h27,8'h27,8'h27,8'h20,8'h20,8'h54,8'h30,8'h4a,8'h88,8'hb7,8'hc6,8'hc6,8'hc5,8'hc1,8'hbb,8'h9c,8'h5d,8'h35,8'h2e,8'h8e,8'hb6,8'hb4,8'hb2,8'hb4,8'had,8'h96,8'h4e,8'h6f,8'h3a,8'h00,8'h2b,8'h3e,8'h26,8'h2c,8'h22,8'h00,8'h4f,8'h47,8'h4d,8'h91,8'h95,8'h93,8'h94,8'h79,8'h34,8'h45,8'h32,8'h00,8'h00,8'h00,8'h00,8'h3a,8'h48,8'h40,8'h81,8'h88,8'h87,8'h86,8'h84,8'h86,8'h79,8'h42,8'h59,8'h3d,8'h00,8'h21,8'h23,8'h25,8'h24,8'h26,8'h2b,8'h2d,8'h34,8'h34,8'h4c,8'h31,8'h0a,8'h00,8'h41,8'h6e,8'h36,8'h15,8'h24,8'h51,8'h68,8'h62,8'h5e,8'h5f,8'h5a,8'h54,8'h4a,8'h2c,8'h21,8'h4b,8'h58,8'h56,8'h57,8'h57,8'h55,8'h3c,8'h41,8'h8e,8'h2a,8'h1f,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h27,8'h25,8'h00,8'h2d,8'h79,8'h37,8'h5f,8'ha6,8'ha9,8'ha8,8'ha6,8'ha5,8'ha7,8'ha6,8'h9c,8'h4c,8'h6a,8'h6a,8'h00,8'h1f,8'h31,8'h45,8'h43,8'h23,8'h25,8'h24,8'h24,8'h25,8'h24,8'h25,8'h24,8'h23,8'h24,8'h24,8'h2b,8'h43,8'h3f,8'h2d,8'h23,8'h20,8'h00,8'h00,8'h33,8'h4e,8'h35,8'h7a,8'h93,8'h8c,8'h8a,8'h89,8'h8a,8'h72,8'h33,8'h67,8'h6e,8'h00,8'h2b,8'h3f,8'h1c,8'h00,8'h44,8'h47,8'h36,8'h79,8'h81,8'h83,8'h81,8'h7f,8'h80,8'h7f,8'h72,8'h69,8'h5e,8'h46,8'h2f,8'h3e,8'h77,8'h7b,8'h79,8'h78,8'h77,8'h75,8'h45,8'h4e,8'h63,8'h00,8'h2e,8'h3d,8'h30,8'h2a,8'h23,8'h00,8'h00,8'h3e,8'h37,8'h63,8'h6b,8'h6e,8'h6d,8'h6b,8'h6d,8'h64,8'h4a,8'h38,8'h6d,8'h20,8'h24,8'h27,8'h27,8'h27,8'h07,8'h30,8'h3c,8'h27,8'h4a,8'h5e,8'h60,8'h5f,8'h5b,8'h50,8'h39,8'h3f,8'h49,8'h47,8'h57,8'h32,8'h3d,8'h48,8'h49,8'h48,8'h47,8'h43,8'h36,8'h2b,8'h70,8'h2b,8'h00,8'h50,8'h48,8'h29,8'h2c,8'h22,8'h00,8'h60,8'h33,8'h28,8'h3d,8'h40,8'h41,8'h41,8'h27,8'h32,8'h4e,8'h00,8'h00,8'h10,8'h07,8'h00,8'h4b,8'h30,8'h2b,8'h3a,8'h41,8'h42,8'h44,8'h41,8'h3b,8'h28,8'h2d,8'h64,8'h23,8'h01,8'h1f,8'h24,8'h25,8'h25,8'h31,8'h36,8'h2f,8'h32,8'h2b,8'h36,8'h2c,8'h00,8'h00,8'h57,8'h3e,8'h2c,8'h3e,8'h44,8'h47,8'h47,8'h43,8'h3e,8'h2a,8'h24,8'h33,8'h44,8'h51,8'h28,8'h3d,8'h44,8'h46,8'h49,8'h47,8'h3f,8'h29,8'h43,8'h8b,8'h29,8'h20,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h22,8'h00,8'h61,8'h64,8'h24,8'h36,8'h45,8'h48,8'h4c,8'h4d,8'h4d,8'h51,8'h4f,8'h43,8'h2c,8'h74,8'h5d,8'h00,8'h3e,8'h40,8'h27,8'h23,8'h23,8'h24,8'h25,8'h26,8'h24,8'h25,8'h26,8'h24,8'h24,8'h28,8'h33,8'h4c,8'h54,8'h50,8'h32,8'h21,8'h00,8'h00,8'h2e,8'h52,8'h31,8'h44,8'h59,8'h5f,8'h5d,8'h61,8'h5f,8'h59,8'h52,8'h3d,8'h3f,8'h80,8'h3c,8'h00,8'h20,8'h00,8'h00,8'h4e,8'h41,8'h38,8'h50,8'h53,8'h5e,8'h5c,8'h59,8'h54,8'h39,8'h2a,8'h4f,8'h65,8'h68,8'h47,8'h37,8'h5a,8'h62,8'h64,8'h64,8'h5f,8'h56,8'h32,8'h53,8'h61,8'h00,8'h44,8'h37,8'h22,8'h2d,8'h27,8'h00,8'h00,8'h41,8'h38,8'h61,8'h6b,8'h73,8'h70,8'h6f,8'h6c,8'h65,8'h47,8'h37,8'h70,8'h21,8'h24,8'h27,8'h27,8'h26,8'h00,8'h44,8'h34,8'h4e,8'h68,8'h6d,8'h6f,8'h75,8'h6c,8'h46,8'h2e,8'h59,8'h62,8'h37,8'h32,8'h30,8'h59,8'h7a,8'h7a,8'h77,8'h77,8'h70,8'h55,8'h40,8'h76,8'h26,8'h00,8'h47,8'h47,8'h2e,8'h27,8'h15,8'h1c,8'h63,8'h2f,8'h53,8'h6f,8'h75,8'h77,8'h6f,8'h37,8'h47,8'h4e,8'h00,8'h00,8'h26,8'h32,8'h47,8'h38,8'h2c,8'h60,8'h77,8'h7b,8'h7c,8'h77,8'h6f,8'h61,8'h38,8'h4d,8'h56,8'h00,8'h0d,8'h21,8'h23,8'h24,8'h26,8'h28,8'h27,8'h2a,8'h2a,8'h25,8'h42,8'h32,8'h00,8'h24,8'h47,8'h32,8'h5a,8'h6c,8'h72,8'h72,8'h70,8'h61,8'h41,8'h3d,8'h59,8'h54,8'h25,8'h3a,8'h2f,8'h60,8'h72,8'h7a,8'h78,8'h73,8'h66,8'h3a,8'h46,8'h8b,8'h27,8'h1e,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h00,8'h00},
'{8'h00,8'h00,8'h27,8'h26,8'h12,8'h27,8'h7d,8'h44,8'h2e,8'h4e,8'h5c,8'h61,8'h66,8'h6d,8'h71,8'h71,8'h6e,8'h54,8'h31,8'h71,8'h59,8'h00,8'h24,8'h28,8'h24,8'h24,8'h25,8'h25,8'h26,8'h24,8'h24,8'h24,8'h36,8'h3f,8'h2a,8'h33,8'h39,8'h53,8'h30,8'h35,8'h20,8'h00,8'h00,8'h31,8'h52,8'h32,8'h45,8'h70,8'h80,8'h81,8'h84,8'h82,8'h81,8'h7c,8'h77,8'h61,8'h30,8'h6a,8'h63,8'h00,8'h00,8'h00,8'h00,8'h58,8'h3c,8'h4e,8'h6e,8'h74,8'h7a,8'h79,8'h74,8'h55,8'h34,8'h5c,8'h5f,8'h26,8'h2e,8'h39,8'h48,8'h72,8'h7e,8'h82,8'h81,8'h77,8'h6b,8'h3e,8'h58,8'h59,8'h00,8'h41,8'h3b,8'h2b,8'h30,8'h23,8'h00,8'h00,8'h3e,8'h41,8'h6e,8'h7f,8'h83,8'h83,8'h80,8'h7e,8'h76,8'h54,8'h39,8'h6f,8'h20,8'h24,8'h27,8'h27,8'h23,8'h00,8'h4b,8'h34,8'h5c,8'h75,8'h7b,8'h7e,8'h7c,8'h6c,8'h3e,8'h5b,8'h4d,8'h00,8'h00,8'h26,8'h36,8'h65,8'h84,8'h86,8'h84,8'h83,8'h7d,8'h61,8'h44,8'h79,8'h1e,8'h07,8'h2e,8'h4f,8'h37,8'h23,8'h00,8'h33,8'h5e,8'h2f,8'h63,8'h7b,8'h81,8'h84,8'h7b,8'h36,8'h55,8'h6f,8'h38,8'h45,8'h50,8'h45,8'h2f,8'h2f,8'h54,8'h79,8'h7f,8'h81,8'h7e,8'h78,8'h68,8'h47,8'h30,8'h62,8'h2a,8'h00,8'h35,8'h26,8'h24,8'h25,8'h29,8'h2c,8'h24,8'h28,8'h48,8'h28,8'h26,8'h21,8'h00,8'h2f,8'h41,8'h38,8'h66,8'h74,8'h7a,8'h78,8'h71,8'h4b,8'h3b,8'h54,8'h36,8'h00,8'h00,8'h34,8'h31,8'h66,8'h79,8'h7f,8'h7b,8'h72,8'h67,8'h3b,8'h4e,8'h8b,8'h1f,8'h15,8'h27,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h26,8'h24,8'h22,8'h26,8'h27,8'h00},
'{8'h00,8'h00,8'h27,8'h25,8'h00,8'h4e,8'h7a,8'h2d,8'h42,8'h5b,8'h66,8'h70,8'h7a,8'h82,8'h84,8'h7f,8'h7a,8'h62,8'h35,8'h67,8'h6a,8'h00,8'h01,8'h21,8'h23,8'h23,8'h24,8'h24,8'h26,8'h25,8'h24,8'h24,8'h37,8'h49,8'h33,8'h3c,8'h2c,8'h28,8'h1c,8'h00,8'h00,8'h17,8'h42,8'h4a,8'h46,8'h55,8'h74,8'h81,8'h8b,8'h8b,8'h89,8'h88,8'h87,8'h84,8'h80,8'h73,8'h44,8'h45,8'h7b,8'h2c,8'h00,8'h00,8'h00,8'h56,8'h34,8'h59,8'h75,8'h7a,8'h7f,8'h7e,8'h6f,8'h45,8'h4f,8'h4f,8'h00,8'h00,8'h27,8'h32,8'h50,8'h75,8'h81,8'h85,8'h84,8'h7d,8'h6b,8'h35,8'h5c,8'h5c,8'h00,8'h3c,8'h2a,8'h23,8'h22,8'h04,8'h00,8'h00,8'h40,8'h40,8'h6c,8'h7d,8'h81,8'h81,8'h81,8'h80,8'h75,8'h56,8'h3b,8'h6e,8'h1d,8'h24,8'h27,8'h27,8'h22,8'h20,8'h4d,8'h39,8'h68,8'h76,8'h7b,8'h7e,8'h7a,8'h5e,8'h44,8'h60,8'h00,8'h00,8'h00,8'h2e,8'h3f,8'h69,8'h82,8'h84,8'h84,8'h82,8'h7f,8'h5b,8'h45,8'h76,8'h00,8'h00,8'h22,8'h32,8'h2a,8'h01,8'h00,8'h4a,8'h4d,8'h33,8'h67,8'h7c,8'h83,8'h86,8'h7f,8'h36,8'h3c,8'h5e,8'h4b,8'h46,8'h46,8'h45,8'h4f,8'h67,8'h77,8'h7d,8'h7b,8'h74,8'h65,8'h4d,8'h43,8'h46,8'h50,8'h42,8'h00,8'h22,8'h4a,8'h38,8'h2b,8'h26,8'h26,8'h28,8'h28,8'h2b,8'h3a,8'h2b,8'h26,8'h0c,8'h00,8'h38,8'h3e,8'h46,8'h6d,8'h7b,8'h80,8'h7c,8'h6d,8'h41,8'h51,8'h32,8'h00,8'h00,8'h00,8'h38,8'h35,8'h68,8'h7a,8'h7d,8'h7b,8'h71,8'h66,8'h38,8'h53,8'h89,8'h20,8'h1c,8'h26,8'h00,8'h26,8'h25,8'h25,8'h25,8'h22,8'h0c,8'h00,8'h08,8'h28,8'h27,8'h27},
'{8'h00,8'h27,8'h27,8'h22,8'h00,8'h72,8'h5e,8'h2b,8'h52,8'h61,8'h6e,8'h79,8'h85,8'h8d,8'h8a,8'h85,8'h81,8'h6f,8'h40,8'h55,8'h80,8'h12,8'h00,8'h1c,8'h23,8'h22,8'h24,8'h23,8'h24,8'h24,8'h24,8'h27,8'h2d,8'h25,8'h2d,8'h34,8'h21,8'h00,8'h00,8'h00,8'h31,8'h51,8'h4a,8'h4b,8'h67,8'h7c,8'h87,8'h8b,8'h8e,8'h8f,8'h91,8'h8d,8'h8b,8'h8a,8'h86,8'h7b,8'h60,8'h2f,8'h6c,8'h60,8'h00,8'h00,8'h20,8'h52,8'h34,8'h64,8'h7a,8'h80,8'h83,8'h7f,8'h66,8'h44,8'h62,8'h14,8'h18,8'h19,8'h30,8'h35,8'h5b,8'h79,8'h88,8'h89,8'h86,8'h80,8'h6e,8'h33,8'h61,8'h63,8'h00,8'h19,8'h15,8'h00,8'h00,8'h00,8'h00,8'h43,8'h4a,8'h42,8'h6d,8'h7c,8'h85,8'h86,8'h87,8'h83,8'h78,8'h56,8'h3d,8'h6e,8'h19,8'h24,8'h27,8'h27,8'h1b,8'h2f,8'h48,8'h41,8'h70,8'h78,8'h7e,8'h7e,8'h7b,8'h53,8'h54,8'h57,8'h00,8'h24,8'h00,8'h33,8'h43,8'h70,8'h85,8'h88,8'h86,8'h82,8'h7c,8'h50,8'h42,8'h72,8'h00,8'h03,8'h1e,8'h15,8'h00,8'h00,8'h00,8'h5b,8'h3d,8'h40,8'h6e,8'h7d,8'h86,8'h88,8'h86,8'h51,8'h39,8'h47,8'h4f,8'h63,8'h72,8'h73,8'h79,8'h7d,8'h7b,8'h75,8'h68,8'h4c,8'h30,8'h36,8'h54,8'h5a,8'h24,8'h00,8'h01,8'h27,8'h2e,8'h55,8'h40,8'h23,8'h24,8'h25,8'h31,8'h46,8'h3b,8'h44,8'h31,8'h00,8'h00,8'h45,8'h39,8'h51,8'h75,8'h7f,8'h81,8'h7e,8'h68,8'h42,8'h5d,8'h23,8'h21,8'h20,8'h00,8'h36,8'h37,8'h6b,8'h7d,8'h7d,8'h7a,8'h70,8'h67,8'h37,8'h58,8'h8a,8'h1d,8'h0f,8'h23,8'h21,8'h1d,8'h01,8'h1f,8'h32,8'h32,8'h00,8'h00,8'h23,8'h29,8'h27,8'h00},
'{8'h00,8'h27,8'h26,8'h09,8'h1b,8'h82,8'h41,8'h33,8'h58,8'h67,8'h7a,8'h81,8'h87,8'h90,8'h8d,8'h8d,8'h89,8'h79,8'h4a,8'h3d,8'h7f,8'h47,8'h00,8'h00,8'h1f,8'h21,8'h21,8'h22,8'h23,8'h24,8'h23,8'h22,8'h22,8'h23,8'h1e,8'h03,8'h00,8'h00,8'h13,8'h4c,8'h52,8'h44,8'h5d,8'h70,8'h7d,8'h85,8'h8c,8'h8f,8'h8f,8'h90,8'h93,8'h8f,8'h8d,8'h8b,8'h86,8'h7d,8'h6f,8'h3c,8'h4c,8'h7a,8'h1f,8'h00,8'h2d,8'h51,8'h37,8'h68,8'h7e,8'h86,8'h86,8'h7b,8'h61,8'h43,8'h5c,8'h01,8'h23,8'h14,8'h32,8'h32,8'h65,8'h7f,8'h8a,8'h89,8'h87,8'h83,8'h72,8'h33,8'h5f,8'h62,8'h00,8'h00,8'h00,8'h00,8'h01,8'h40,8'h68,8'h8c,8'h51,8'h43,8'h71,8'h84,8'h8a,8'h88,8'h88,8'h81,8'h78,8'h56,8'h3b,8'h6f,8'h10,8'h24,8'h27,8'h27,8'h12,8'h41,8'h44,8'h4d,8'h79,8'h7f,8'h7f,8'h80,8'h7a,8'h4b,8'h60,8'h52,8'h00,8'h1a,8'h00,8'h38,8'h42,8'h72,8'h86,8'h8a,8'h8d,8'h89,8'h7f,8'h4d,8'h42,8'h6d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h70,8'h36,8'h4d,8'h78,8'h81,8'h89,8'h8c,8'h89,8'h80,8'h7d,8'h7d,8'h7c,8'h7d,8'h81,8'h80,8'h7d,8'h7c,8'h6f,8'h56,8'h42,8'h35,8'h4b,8'h5d,8'h3d,8'h00,8'h00,8'h0b,8'h24,8'h22,8'h26,8'h2f,8'h29,8'h24,8'h24,8'h23,8'h2c,8'h40,8'h4a,8'h6d,8'h42,8'h00,8'h00,8'h48,8'h3a,8'h59,8'h78,8'h7e,8'h81,8'h7c,8'h61,8'h42,8'h5b,8'h0a,8'h06,8'h01,8'h36,8'h36,8'h3e,8'h72,8'h80,8'h7e,8'h7b,8'h75,8'h68,8'h36,8'h56,8'h85,8'h00,8'h00,8'h13,8'h08,8'h2f,8'h57,8'h82,8'h9e,8'h66,8'h19,8'h1a,8'h27,8'h00,8'h00,8'h00},
'{8'h00,8'h26,8'h22,8'h00,8'h46,8'h85,8'h2f,8'h44,8'h61,8'h6f,8'h7e,8'h85,8'h8c,8'h8f,8'h91,8'h92,8'h8e,8'h84,8'h6a,8'h3b,8'h4e,8'h7a,8'h40,8'h00,8'h00,8'h00,8'h00,8'h02,8'h09,8'h09,8'h05,8'h00,8'h00,8'h00,8'h00,8'h02,8'h44,8'h55,8'h49,8'h4a,8'h52,8'h67,8'h7a,8'h83,8'h87,8'h8c,8'h90,8'h91,8'h91,8'h8f,8'h93,8'h8e,8'h8b,8'h8a,8'h85,8'h80,8'h78,8'h5a,8'h36,8'h73,8'h50,8'h00,8'h46,8'h4a,8'h3e,8'h6e,8'h7f,8'h85,8'h86,8'h7b,8'h5a,8'h43,8'h55,8'h00,8'h00,8'h00,8'h3f,8'h32,8'h6b,8'h84,8'h8b,8'h8a,8'h89,8'h83,8'h71,8'h32,8'h5c,8'h57,8'h00,8'h00,8'h3e,8'h69,8'h76,8'h6a,8'h71,8'h9f,8'h4e,8'h41,8'h70,8'h81,8'h87,8'h87,8'h86,8'h82,8'h78,8'h58,8'h3f,8'h72,8'h0b,8'h23,8'h27,8'h26,8'h1d,8'h4b,8'h36,8'h5b,8'h7b,8'h82,8'h82,8'h83,8'h77,8'h43,8'h6a,8'h40,8'h00,8'h2b,8'h4a,8'h37,8'h50,8'h7e,8'h89,8'h8b,8'h8e,8'h8b,8'h80,8'h4d,8'h46,8'h6f,8'h00,8'h00,8'h00,8'h05,8'h49,8'h57,8'h61,8'h77,8'h2f,8'h5d,8'h7d,8'h82,8'h85,8'h87,8'h88,8'h84,8'h83,8'h7f,8'h7f,8'h80,8'h84,8'h82,8'h7b,8'h69,8'h44,8'h47,8'h53,8'h3e,8'h2e,8'h0e,8'h00,8'h05,8'h26,8'h2c,8'h2b,8'h24,8'h24,8'h24,8'h24,8'h24,8'h24,8'h29,8'h41,8'h4b,8'h4d,8'h49,8'h33,8'h00,8'h00,8'h4b,8'h38,8'h64,8'h7b,8'h82,8'h83,8'h78,8'h5a,8'h46,8'h57,8'h00,8'h21,8'h56,8'h56,8'h2e,8'h4d,8'h75,8'h7f,8'h7b,8'h7a,8'h79,8'h6a,8'h34,8'h56,8'h90,8'h3f,8'h47,8'h70,8'h75,8'h64,8'h72,8'hae,8'h74,8'h2a,8'h20,8'h27,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h26,8'h12,8'h00,8'h63,8'h74,8'h2a,8'h4e,8'h65,8'h76,8'h82,8'h89,8'h8f,8'h90,8'h94,8'h95,8'h92,8'h8b,8'h80,8'h5c,8'h29,8'h49,8'h76,8'h53,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2f,8'h56,8'h68,8'h5a,8'h3e,8'h41,8'h5a,8'h74,8'h82,8'h88,8'h8e,8'h91,8'h90,8'h94,8'h95,8'h92,8'h8e,8'h91,8'h8e,8'h8e,8'h8a,8'h85,8'h84,8'h7c,8'h6b,8'h3f,8'h54,8'h79,8'h20,8'h52,8'h44,8'h43,8'h71,8'h7e,8'h86,8'h84,8'h7b,8'h55,8'h49,8'h53,8'h00,8'h00,8'h49,8'h46,8'h44,8'h74,8'h86,8'h8d,8'h8b,8'h8b,8'h83,8'h6f,8'h2e,8'h5e,8'h67,8'h4a,8'h78,8'h8a,8'h73,8'h43,8'h3c,8'h73,8'h90,8'h4d,8'h44,8'h72,8'h81,8'h86,8'h86,8'h85,8'h81,8'h7a,8'h57,8'h3f,8'h70,8'h06,8'h23,8'h27,8'h25,8'h23,8'h4f,8'h32,8'h64,8'h7d,8'h82,8'h85,8'h83,8'h75,8'h43,8'h7e,8'h5b,8'h52,8'h69,8'h41,8'h3b,8'h6d,8'h86,8'h8c,8'h8c,8'h8c,8'h88,8'h7f,8'h4f,8'h47,8'h88,8'h2f,8'h23,8'h56,8'h6a,8'h54,8'h31,8'h4d,8'h6d,8'h29,8'h5a,8'h78,8'h7f,8'h80,8'h83,8'h82,8'h82,8'h82,8'h7c,8'h7b,8'h7b,8'h82,8'h80,8'h72,8'h43,8'h40,8'h5d,8'h27,8'h00,8'h00,8'h00,8'h1e,8'h3d,8'h52,8'h34,8'h34,8'h2b,8'h24,8'h24,8'h22,8'h24,8'h24,8'h2b,8'h50,8'h5d,8'h5e,8'h4b,8'h22,8'h00,8'h22,8'h48,8'h39,8'h6a,8'h7d,8'h87,8'h84,8'h7d,8'h56,8'h4d,8'h73,8'h5c,8'h73,8'h56,8'h2d,8'h41,8'h63,8'h72,8'h7c,8'h7c,8'h7d,8'h78,8'h67,8'h35,8'h5a,8'hae,8'h99,8'h8c,8'h6d,8'h44,8'h29,8'h5d,8'h69,8'h08,8'h13,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00},
'{8'h27,8'h26,8'h07,8'h00,8'h73,8'h5a,8'h2f,8'h55,8'h65,8'h75,8'h84,8'h8b,8'h8f,8'h93,8'h97,8'h93,8'h91,8'h8f,8'h89,8'h7a,8'h53,8'h2e,8'h41,8'h63,8'h61,8'h50,8'h48,8'h38,8'h33,8'h3c,8'h3f,8'h4a,8'h65,8'h72,8'h63,8'h47,8'h3a,8'h57,8'h6f,8'h7f,8'h87,8'h8d,8'h91,8'h92,8'h91,8'h90,8'h8f,8'h92,8'h91,8'h91,8'h8f,8'h8d,8'h8e,8'h8b,8'h86,8'h84,8'h7e,8'h76,8'h50,8'h3a,8'h7b,8'h5f,8'h64,8'h3f,8'h4c,8'h7a,8'h84,8'h88,8'h8a,8'h83,8'h57,8'h49,8'h6b,8'h4d,8'h65,8'h60,8'h42,8'h60,8'h7f,8'h89,8'h8b,8'h8b,8'h8b,8'h84,8'h76,8'h35,8'h50,8'h86,8'h82,8'h71,8'h45,8'h22,8'h2c,8'h64,8'h61,8'h4a,8'h41,8'h47,8'h78,8'h83,8'h86,8'h87,8'h84,8'h81,8'h78,8'h54,8'h41,8'h6f,8'h05,8'h23,8'h27,8'h23,8'h25,8'h43,8'h36,8'h69,8'h7d,8'h83,8'h88,8'h86,8'h75,8'h42,8'h7a,8'h7d,8'h5f,8'h3d,8'h3e,8'h69,8'h80,8'h86,8'h89,8'h8c,8'h8b,8'h89,8'h80,8'h55,8'h41,8'h8e,8'h76,8'h6a,8'h57,8'h2d,8'h1a,8'h33,8'h77,8'h6a,8'h2a,8'h60,8'h75,8'h7c,8'h79,8'h7a,8'h7a,8'h7a,8'h6d,8'h5f,8'h55,8'h4b,8'h5b,8'h73,8'h5a,8'h35,8'h5f,8'h2b,8'h00,8'h00,8'h11,8'h23,8'h32,8'h4a,8'h55,8'h40,8'h4e,8'h25,8'h23,8'h28,8'h30,8'h2a,8'h24,8'h24,8'h29,8'h49,8'h4a,8'h4a,8'h1d,8'h00,8'h2f,8'h44,8'h42,8'h72,8'h80,8'h87,8'h83,8'h7d,8'h50,8'h4a,8'h87,8'h73,8'h47,8'h32,8'h47,8'h65,8'h74,8'h7a,8'h7c,8'h7f,8'h80,8'h7e,8'h6a,8'h34,8'h49,8'h81,8'h60,8'h3c,8'h18,8'h1d,8'h4e,8'h6c,8'h26,8'h17,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h27,8'h26,8'h00,8'h0e,8'h78,8'h48,8'h38,8'h59,8'h6a,8'h7a,8'h83,8'h89,8'h8f,8'h91,8'h97,8'h98,8'h94,8'h90,8'h8c,8'h87,8'h80,8'h72,8'h59,8'h48,8'h44,8'h45,8'h49,8'h45,8'h45,8'h4a,8'h44,8'h40,8'h46,8'h4e,8'h53,8'h61,8'h71,8'h81,8'h83,8'h8b,8'h8f,8'h91,8'h91,8'h92,8'h90,8'h91,8'h8f,8'h92,8'h90,8'h8f,8'h91,8'h8e,8'h8b,8'h8c,8'h88,8'h82,8'h7c,8'h75,8'h64,8'h33,8'h55,8'h96,8'h73,8'h2e,8'h58,8'h7c,8'h84,8'h8b,8'h8b,8'h88,8'h67,8'h3d,8'h45,8'h42,8'h4f,8'h58,8'h6b,8'h7a,8'h84,8'h8b,8'h8a,8'h8b,8'h8b,8'h83,8'h7b,8'h54,8'h2f,8'h36,8'h3f,8'h39,8'h25,8'h43,8'h73,8'h45,8'h00,8'h34,8'h3e,8'h48,8'h78,8'h83,8'h86,8'h86,8'h84,8'h81,8'h76,8'h52,8'h42,8'h72,8'h09,8'h24,8'h27,8'h23,8'h3b,8'h40,8'h48,8'h74,8'h81,8'h88,8'h87,8'h88,8'h80,8'h4a,8'h3c,8'h4a,8'h58,8'h68,8'h75,8'h80,8'h84,8'h88,8'h8d,8'h90,8'h8b,8'h89,8'h83,8'h64,8'h29,8'h36,8'h39,8'h32,8'h2c,8'h23,8'h46,8'h51,8'h6a,8'h58,8'h30,8'h61,8'h6c,8'h72,8'h6d,8'h63,8'h55,8'h46,8'h3d,8'h45,8'h5a,8'h3a,8'h30,8'h61,8'h40,8'h54,8'h4d,8'h00,8'h00,8'h0d,8'h1c,8'h18,8'h1a,8'h19,8'h1b,8'h20,8'h26,8'h15,8'h1c,8'h2d,8'h67,8'h43,8'h2c,8'h3c,8'h35,8'h2b,8'h24,8'h25,8'h05,8'h00,8'h42,8'h3c,8'h4c,8'h76,8'h80,8'h88,8'h85,8'h7e,8'h5a,8'h2a,8'h38,8'h46,8'h53,8'h64,8'h6f,8'h78,8'h7a,8'h7d,8'h7e,8'h7e,8'h7f,8'h7c,8'h6d,8'h44,8'h27,8'h2f,8'h32,8'h28,8'h20,8'h56,8'h63,8'h2c,8'h1f,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h27,8'h25,8'h00,8'h26,8'h7c,8'h3a,8'h41,8'h5c,8'h6d,8'h80,8'h85,8'h88,8'h8e,8'h92,8'h93,8'h95,8'h97,8'h93,8'h91,8'h8e,8'h8a,8'h85,8'h7c,8'h6d,8'h62,8'h57,8'h4b,8'h46,8'h47,8'h4a,8'h4d,8'h59,8'h64,8'h6c,8'h74,8'h7f,8'h85,8'h87,8'h8d,8'h90,8'h90,8'h91,8'h93,8'h93,8'h8f,8'h93,8'h91,8'h92,8'h90,8'h91,8'h91,8'h8d,8'h86,8'h86,8'h82,8'h7f,8'h7b,8'h71,8'h64,8'h38,8'h34,8'h8d,8'h69,8'h2b,8'h5f,8'h7e,8'h85,8'h8c,8'h8a,8'h88,8'h80,8'h62,8'h55,8'h61,8'h72,8'h77,8'h7e,8'h82,8'h85,8'h8a,8'h88,8'h87,8'h86,8'h80,8'h7d,8'h71,8'h52,8'h4c,8'h4b,8'h30,8'h45,8'h7b,8'h4c,8'h00,8'h00,8'h3a,8'h3e,8'h4a,8'h75,8'h7f,8'h81,8'h83,8'h80,8'h7d,8'h77,8'h52,8'h3f,8'h72,8'h06,8'h23,8'h27,8'h1e,8'h42,8'h3a,8'h50,8'h78,8'h81,8'h86,8'h85,8'h89,8'h89,8'h79,8'h6e,8'h77,8'h7d,8'h82,8'h80,8'h80,8'h85,8'h88,8'h8e,8'h8e,8'h8b,8'h89,8'h83,8'h77,8'h4e,8'h39,8'h40,8'h39,8'h2e,8'h56,8'h57,8'h00,8'h5a,8'h4e,8'h31,8'h5b,8'h5f,8'h55,8'h44,8'h33,8'h33,8'h49,8'h53,8'h5f,8'h83,8'h45,8'h3a,8'h55,8'h3c,8'h6a,8'h21,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2f,8'h27,8'h4c,8'h64,8'h42,8'h2a,8'h23,8'h23,8'h00,8'h00,8'h50,8'h32,8'h54,8'h7a,8'h82,8'h86,8'h88,8'h86,8'h78,8'h59,8'h5a,8'h6a,8'h77,8'h79,8'h7b,8'h7c,8'h77,8'h7a,8'h7c,8'h79,8'h76,8'h77,8'h6e,8'h60,8'h4a,8'h44,8'h3b,8'h27,8'h54,8'h61,8'h22,8'h11,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h27,8'h26,8'h00,8'h2c,8'h80,8'h36,8'h41,8'h5c,8'h6b,8'h7d,8'h85,8'h8a,8'h8e,8'h90,8'h95,8'h97,8'h93,8'h92,8'h92,8'h90,8'h8d,8'h8a,8'h87,8'h81,8'h80,8'h7b,8'h72,8'h71,8'h73,8'h72,8'h74,8'h7d,8'h80,8'h7f,8'h7f,8'h86,8'h8a,8'h89,8'h90,8'h94,8'h94,8'h98,8'h95,8'h91,8'h91,8'h92,8'h90,8'h8f,8'h8d,8'h8d,8'h8d,8'h86,8'h82,8'h7e,8'h79,8'h73,8'h65,8'h4d,8'h42,8'h45,8'h65,8'h9d,8'h5f,8'h32,8'h66,8'h7f,8'h87,8'h8c,8'h8a,8'h88,8'h89,8'h85,8'h83,8'h83,8'h85,8'h82,8'h82,8'h82,8'h82,8'h83,8'h84,8'h85,8'h85,8'h84,8'h7d,8'h73,8'h67,8'h57,8'h45,8'h55,8'h77,8'h48,8'h00,8'h00,8'h00,8'h3d,8'h3f,8'h4c,8'h75,8'h7f,8'h82,8'h82,8'h82,8'h7e,8'h78,8'h4c,8'h3c,8'h6f,8'h11,8'h24,8'h26,8'h1b,8'h44,8'h35,8'h60,8'h7a,8'h81,8'h86,8'h86,8'h8a,8'h8a,8'h8a,8'h8c,8'h88,8'h86,8'h84,8'h81,8'h82,8'h85,8'h85,8'h87,8'h86,8'h85,8'h81,8'h81,8'h7c,8'h71,8'h63,8'h4b,8'h3f,8'h56,8'h58,8'h00,8'h00,8'h6a,8'h59,8'h27,8'h40,8'h45,8'h4d,8'h48,8'h45,8'h53,8'h4f,8'h24,8'h4d,8'h57,8'h38,8'h57,8'h47,8'h4c,8'h61,8'h00,8'h01,8'h24,8'h33,8'h3f,8'h3e,8'h3f,8'h41,8'h42,8'h41,8'h41,8'h42,8'h2b,8'h00,8'h00,8'h00,8'h14,8'h2c,8'h2d,8'h24,8'h24,8'h23,8'h00,8'h00,8'h59,8'h2f,8'h5d,8'h7d,8'h82,8'h85,8'h86,8'h87,8'h88,8'h83,8'h80,8'h7d,8'h7d,8'h7a,8'h77,8'h77,8'h74,8'h70,8'h6c,8'h70,8'h72,8'h70,8'h67,8'h61,8'h54,8'h3c,8'h2d,8'h56,8'h6b,8'h27,8'h1b,8'h29,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h27,8'h25,8'h00,8'h2c,8'h81,8'h34,8'h3f,8'h5e,8'h6a,8'h7b,8'h86,8'h8b,8'h8d,8'h8f,8'h92,8'h92,8'h94,8'h94,8'h91,8'h8f,8'h8f,8'h8d,8'h8f,8'h8d,8'h8b,8'h86,8'h80,8'h83,8'h86,8'h88,8'h88,8'h85,8'h84,8'h83,8'h83,8'h86,8'h7b,8'h69,8'h86,8'h92,8'h97,8'h99,8'h94,8'h8f,8'h8d,8'h8e,8'h8c,8'h8c,8'h8b,8'h88,8'h84,8'h7d,8'h7a,8'h74,8'h62,8'h4b,8'h35,8'h40,8'h6d,8'h8d,8'h72,8'h78,8'h4d,8'h36,8'h6e,8'h81,8'h88,8'h89,8'h89,8'h8c,8'h8a,8'h85,8'h88,8'h87,8'h80,8'h7f,8'h7d,8'h7c,8'h75,8'h70,8'h7f,8'h80,8'h80,8'h7e,8'h74,8'h6d,8'h53,8'h3f,8'h70,8'h88,8'h39,8'h00,8'h23,8'h26,8'h00,8'h3d,8'h3f,8'h4e,8'h75,8'h7e,8'h82,8'h7f,8'h7f,8'h7e,8'h6f,8'h3e,8'h49,8'h7e,8'h13,8'h24,8'h23,8'h1b,8'h4c,8'h3c,8'h68,8'h7d,8'h85,8'h86,8'h89,8'h8b,8'h89,8'h88,8'h88,8'h87,8'h86,8'h83,8'h7f,8'h7d,8'h78,8'h77,8'h7f,8'h80,8'h82,8'h82,8'h7d,8'h76,8'h67,8'h47,8'h46,8'h6e,8'h4c,8'h00,8'h00,8'h00,8'h58,8'h83,8'h60,8'h64,8'h6d,8'h62,8'h45,8'h1a,8'h00,8'h00,8'h21,8'h5e,8'h2e,8'h51,8'h66,8'h39,8'h5d,8'h84,8'h72,8'h7b,8'h75,8'h70,8'h66,8'h5c,8'h5a,8'h5a,8'h62,8'h6b,8'h7c,8'h8f,8'h8d,8'h7b,8'h5a,8'h29,8'h00,8'h00,8'h00,8'h18,8'h23,8'h23,8'h00,8'h15,8'h4f,8'h30,8'h64,8'h7c,8'h83,8'h84,8'h83,8'h85,8'h83,8'h80,8'h7d,8'h7d,8'h7a,8'h75,8'h6b,8'h65,8'h54,8'h37,8'h42,8'h67,8'h6a,8'h68,8'h63,8'h56,8'h36,8'h29,8'h63,8'h68,8'h20,8'h1b,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h27,8'h26,8'h00,8'h2c,8'h82,8'h36,8'h3a,8'h58,8'h68,8'h78,8'h83,8'h8c,8'h8e,8'h8f,8'h91,8'h93,8'h93,8'h90,8'h90,8'h8e,8'h8e,8'h90,8'h91,8'h91,8'h8c,8'h88,8'h84,8'h87,8'h86,8'h86,8'h86,8'h84,8'h81,8'h80,8'h7f,8'h6e,8'h43,8'h36,8'h7e,8'h93,8'h92,8'h92,8'h91,8'h8f,8'h8c,8'h8a,8'h84,8'h86,8'h84,8'h80,8'h7b,8'h73,8'h64,8'h4f,8'h3b,8'h41,8'h6a,8'h8b,8'h71,8'h3d,8'h00,8'h52,8'h45,8'h3b,8'h71,8'h80,8'h84,8'h88,8'h88,8'h86,8'h87,8'h83,8'h82,8'h80,8'h7d,8'h78,8'h71,8'h66,8'h47,8'h3e,8'h6a,8'h79,8'h79,8'h74,8'h68,8'h55,8'h45,8'h75,8'h88,8'h38,8'h01,8'h24,8'h27,8'h27,8'h06,8'h42,8'h3f,8'h4e,8'h71,8'h7a,8'h7e,8'h7d,8'h7c,8'h77,8'h5f,8'h31,8'h71,8'h7e,8'h00,8'h23,8'h21,8'h26,8'h49,8'h42,8'h6d,8'h7d,8'h81,8'h82,8'h85,8'h87,8'h87,8'h85,8'h84,8'h82,8'h7e,8'h7a,8'h73,8'h64,8'h47,8'h42,8'h70,8'h80,8'h81,8'h7d,8'h7a,8'h6b,8'h48,8'h45,8'h76,8'h4e,8'h00,8'h1e,8'h22,8'h00,8'h03,8'h49,8'h51,8'h3d,8'h21,8'h00,8'h00,8'h00,8'h00,8'h00,8'h61,8'h45,8'h37,8'h61,8'h64,8'h3f,8'h3e,8'h67,8'h61,8'h4a,8'h34,8'h2d,8'h2d,8'h2c,8'h2c,8'h2d,8'h2c,8'h2a,8'h2c,8'h39,8'h4d,8'h6b,8'h90,8'h8c,8'h5a,8'h16,8'h00,8'h00,8'h0f,8'h19,8'h00,8'h2f,8'h49,8'h36,8'h66,8'h7a,8'h83,8'h83,8'h82,8'h83,8'h7f,8'h7c,8'h77,8'h74,8'h6f,8'h66,8'h54,8'h41,8'h2e,8'h25,8'h30,8'h5e,8'h65,8'h65,8'h5b,8'h40,8'h27,8'h61,8'h73,8'h28,8'h13,8'h29,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h27,8'h26,8'h00,8'h1c,8'h83,8'h48,8'h2f,8'h53,8'h64,8'h75,8'h81,8'h86,8'h8a,8'h8c,8'h8f,8'h91,8'h8f,8'h8d,8'h8d,8'h8e,8'h8f,8'h8e,8'h92,8'h8e,8'h86,8'h87,8'h84,8'h85,8'h80,8'h7e,8'h7f,8'h7d,8'h72,8'h68,8'h4e,8'h40,8'h24,8'h40,8'h82,8'h8e,8'h8f,8'h8e,8'h8b,8'h89,8'h8b,8'h86,8'h7e,8'h7a,8'h72,8'h6c,8'h5c,8'h43,8'h43,8'h67,8'h80,8'h7a,8'h5e,8'h41,8'h00,8'h00,8'h00,8'h5e,8'h3b,8'h47,8'h71,8'h79,8'h7f,8'h86,8'h82,8'h81,8'h80,8'h7f,8'h79,8'h75,8'h70,8'h65,8'h4a,8'h4d,8'h5e,8'h34,8'h55,8'h70,8'h72,8'h64,8'h4a,8'h59,8'h87,8'h79,8'h2e,8'h0c,8'h24,8'h27,8'h27,8'h26,8'h00,8'h46,8'h41,8'h4d,8'h6c,8'h74,8'h7a,8'h77,8'h72,8'h59,8'h3e,8'h64,8'h99,8'h48,8'h0a,8'h25,8'h18,8'h38,8'h4c,8'h47,8'h6d,8'h7d,8'h81,8'h81,8'h7e,8'h7d,8'h7c,8'h79,8'h7b,8'h74,8'h6f,8'h63,8'h47,8'h56,8'h69,8'h31,8'h57,8'h78,8'h78,8'h74,8'h61,8'h43,8'h60,8'h70,8'h44,8'h18,8'h23,8'h27,8'h26,8'h1f,8'h04,8'h00,8'h00,8'h00,8'h11,8'h22,8'h22,8'h19,8'h00,8'h4a,8'h5c,8'h2e,8'h4a,8'h50,8'h44,8'h30,8'h20,8'h1e,8'h22,8'h29,8'h38,8'h47,8'h53,8'h59,8'h5e,8'h62,8'h62,8'h60,8'h55,8'h4a,8'h43,8'h41,8'h44,8'h54,8'h73,8'h82,8'h53,8'h00,8'h00,8'h00,8'h00,8'h43,8'h3f,8'h3e,8'h65,8'h75,8'h7e,8'h7f,8'h7c,8'h78,8'h72,8'h72,8'h6d,8'h66,8'h52,8'h3a,8'h34,8'h58,8'h75,8'h62,8'h2f,8'h51,8'h60,8'h59,8'h39,8'h30,8'h69,8'h64,8'h28,8'h19,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h27,8'h26,8'h09,8'h00,8'h72,8'h5a,8'h28,8'h4f,8'h61,8'h6d,8'h7a,8'h81,8'h84,8'h85,8'h8a,8'h8d,8'h8c,8'h8c,8'h8d,8'h8c,8'h8a,8'h8a,8'h8b,8'h89,8'h87,8'h86,8'h82,8'h80,8'h7c,8'h77,8'h73,8'h6b,8'h56,8'h3a,8'h41,8'h59,8'h30,8'h51,8'h83,8'h8b,8'h8e,8'h89,8'h88,8'h87,8'h85,8'h7f,8'h76,8'h6d,8'h5b,8'h41,8'h36,8'h54,8'h89,8'h99,8'h6c,8'h2b,8'h00,8'h03,8'h22,8'h24,8'h0e,8'h5b,8'h31,8'h49,8'h6d,8'h73,8'h78,8'h7f,8'h7e,8'h7b,8'h79,8'h79,8'h75,8'h66,8'h52,8'h3e,8'h4d,8'h8b,8'h94,8'h41,8'h46,8'h67,8'h64,8'h44,8'h4f,8'h9f,8'h7c,8'h20,8'h0e,8'h27,8'h27,8'h27,8'h27,8'h24,8'h00,8'h51,8'h44,8'h4e,8'h6c,8'h72,8'h71,8'h6a,8'h56,8'h38,8'h67,8'hac,8'h65,8'h00,8'h24,8'h26,8'h0e,8'h48,8'h54,8'h49,8'h6c,8'h79,8'h7a,8'h7b,8'h79,8'h76,8'h73,8'h6f,8'h68,8'h5a,8'h49,8'h42,8'h6b,8'h8f,8'h8b,8'h43,8'h4b,8'h74,8'h73,8'h5f,8'h3a,8'h5f,8'h7d,8'h38,8'h00,8'h26,8'h28,8'h27,8'h00,8'h26,8'h26,8'h26,8'h25,8'h25,8'h26,8'h27,8'h26,8'h16,8'h29,8'h72,8'h2e,8'h27,8'h32,8'h33,8'h38,8'h44,8'h4b,8'h48,8'h3d,8'h2e,8'h29,8'h32,8'h49,8'h60,8'h6a,8'h72,8'h79,8'h7e,8'h7c,8'h7b,8'h74,8'h6c,8'h53,8'h35,8'h2b,8'h65,8'h9b,8'h63,8'h00,8'h00,8'h00,8'h60,8'h3d,8'h3b,8'h63,8'h6d,8'h75,8'h72,8'h71,8'h6d,8'h65,8'h5c,8'h50,8'h3a,8'h29,8'h43,8'h6e,8'h6d,8'h65,8'h74,8'h2d,8'h45,8'h4e,8'h3a,8'h28,8'h6b,8'h72,8'h05,8'h12,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h26,8'h14,8'h00,8'h58,8'h77,8'h2c,8'h44,8'h58,8'h66,8'h75,8'h7c,8'h7e,8'h85,8'h89,8'h8c,8'h8e,8'h8b,8'h8c,8'h89,8'h87,8'h87,8'h86,8'h85,8'h84,8'h81,8'h7b,8'h76,8'h73,8'h6a,8'h59,8'h4a,8'h42,8'h61,8'h93,8'h73,8'h2d,8'h5e,8'h80,8'h87,8'h88,8'h83,8'h80,8'h7c,8'h77,8'h6c,8'h5b,8'h4d,8'h3f,8'h47,8'h7b,8'h99,8'h76,8'h33,8'h00,8'h05,8'h23,8'h27,8'h27,8'h25,8'h0b,8'h65,8'h39,8'h42,8'h68,8'h6f,8'h72,8'h77,8'h74,8'h74,8'h6f,8'h63,8'h58,8'h4a,8'h41,8'h62,8'h89,8'h62,8'h58,8'h4a,8'h3d,8'h52,8'h49,8'h53,8'h92,8'h7c,8'h28,8'h20,8'h27,8'h27,8'h27,8'h27,8'h27,8'h24,8'h00,8'h5b,8'h47,8'h4e,8'h68,8'h6e,8'h65,8'h4b,8'h3c,8'h68,8'hab,8'h70,8'h0b,8'h1c,8'h27,8'h26,8'h09,8'h47,8'h5b,8'h47,8'h66,8'h6d,8'h6f,8'h71,8'h6c,8'h66,8'h60,8'h57,8'h51,8'h44,8'h4d,8'h7a,8'h7a,8'h39,8'h4a,8'h51,8'h42,8'h63,8'h57,8'h45,8'h60,8'h7b,8'h39,8'h1a,8'h25,8'h27,8'h27,8'h00,8'h00,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h24,8'h04,8'h5b,8'h62,8'h2f,8'h3e,8'h58,8'h76,8'h85,8'h7d,8'h77,8'h77,8'h72,8'h75,8'h63,8'h3b,8'h32,8'h40,8'h59,8'h6c,8'h78,8'h7e,8'h83,8'h84,8'h7d,8'h7c,8'h7b,8'h67,8'h47,8'h2d,8'h59,8'h94,8'h61,8'h09,8'h2c,8'h87,8'h56,8'h2f,8'h54,8'h62,8'h69,8'h66,8'h5f,8'h56,8'h45,8'h38,8'h35,8'h3a,8'h63,8'h76,8'h4b,8'h00,8'h2f,8'h6f,8'h2b,8'h39,8'h36,8'h28,8'h5c,8'h79,8'h26,8'h0f,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h27,8'h23,8'h00,8'h30,8'h8f,8'h4a,8'h30,8'h4e,8'h61,8'h6d,8'h75,8'h7d,8'h84,8'h87,8'h87,8'h88,8'h88,8'h87,8'h84,8'h83,8'h82,8'h80,8'h7c,8'h7d,8'h77,8'h6e,8'h65,8'h59,8'h41,8'h41,8'h66,8'h88,8'h8a,8'h87,8'h58,8'h2f,8'h66,8'h7e,8'h84,8'h7d,8'h75,8'h72,8'h69,8'h53,8'h3a,8'h42,8'h6a,8'h89,8'h7e,8'h5b,8'h36,8'h15,8'h21,8'h25,8'h26,8'h27,8'h00,8'h27,8'h24,8'h00,8'h6a,8'h63,8'h2c,8'h4e,8'h60,8'h61,8'h5f,8'h56,8'h49,8'h40,8'h3f,8'h5f,8'h7e,8'h75,8'h54,8'h2e,8'h00,8'h40,8'h5d,8'h26,8'h3a,8'h77,8'h94,8'h59,8'h20,8'h24,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h25,8'h12,8'h63,8'h46,8'h47,8'h61,8'h4c,8'h38,8'h57,8'h95,8'h97,8'h55,8'h20,8'h23,8'h26,8'h27,8'h27,8'h20,8'h36,8'h70,8'h3e,8'h44,8'h4e,8'h4c,8'h49,8'h41,8'h3e,8'h49,8'h69,8'h7f,8'h6e,8'h50,8'h37,8'h11,8'h00,8'h2d,8'h56,8'h34,8'h44,8'h41,8'h74,8'h68,8'h2d,8'h23,8'h28,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h00,8'h2c,8'h86,8'h71,8'h5c,8'h46,8'h39,8'h2c,8'h27,8'h00,8'h00,8'h00,8'h22,8'h73,8'ha0,8'h88,8'h6c,8'h4d,8'h30,8'h4f,8'h6e,8'h77,8'h82,8'h84,8'h85,8'h85,8'h8a,8'h82,8'h76,8'h5b,8'h36,8'h4e,8'h93,8'h85,8'h5e,8'h5c,8'h70,8'h38,8'h2e,8'h41,8'h41,8'h36,8'h2a,8'h30,8'h45,8'h65,8'h6a,8'h54,8'h41,8'h24,8'h02,8'h00,8'h31,8'h81,8'h34,8'h1c,8'h32,8'h6d,8'h66,8'h26,8'h1d,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h27,8'h26,8'h20,8'h00,8'h77,8'h78,8'h29,8'h3f,8'h58,8'h65,8'h6b,8'h76,8'h7b,8'h7f,8'h80,8'h80,8'h81,8'h81,8'h7d,8'h79,8'h79,8'h74,8'h70,8'h6c,8'h65,8'h58,8'h43,8'h33,8'h49,8'h7e,8'h98,8'h78,8'h39,8'h5f,8'h43,8'h3d,8'h6d,8'h76,8'h77,8'h6c,8'h65,8'h55,8'h3a,8'h36,8'h5d,8'h97,8'ha2,8'h69,8'h29,8'h00,8'h15,8'h24,8'h27,8'h27,8'h27,8'h00,8'h00,8'h27,8'h25,8'h01,8'h4a,8'ha1,8'h54,8'h2b,8'h31,8'h2c,8'h2c,8'h34,8'h42,8'h61,8'h84,8'h86,8'h61,8'h33,8'h14,8'h1e,8'h12,8'h39,8'h7a,8'h45,8'h77,8'ha7,8'h57,8'h00,8'h21,8'h27,8'h00,8'h27,8'h27,8'h27,8'h27,8'h27,8'h26,8'h17,8'h66,8'h4b,8'h30,8'h37,8'h2f,8'h66,8'hb1,8'h99,8'h41,8'h00,8'h24,8'h27,8'h27,8'h00,8'h27,8'h26,8'h20,8'h70,8'h76,8'h3e,8'h33,8'h43,8'h52,8'h63,8'h7f,8'h8a,8'h82,8'h5a,8'h2d,8'h00,8'h0c,8'h24,8'h23,8'h21,8'h68,8'h2e,8'h38,8'h79,8'h69,8'h1b,8'h20,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h23,8'h00,8'h1a,8'h4f,8'h3f,8'h24,8'h18,8'h12,8'h0a,8'h0e,8'h00,8'h00,8'h00,8'h4d,8'h9e,8'ha5,8'h62,8'h3b,8'h6f,8'h4d,8'h2e,8'h5e,8'h73,8'h81,8'h85,8'h8b,8'h8a,8'h8a,8'h87,8'h80,8'h76,8'h53,8'h28,8'h6d,8'ha7,8'h43,8'h00,8'h46,8'h68,8'h3e,8'h2a,8'h2b,8'h3d,8'h54,8'h72,8'h74,8'h5e,8'h2c,8'h00,8'h00,8'h22,8'h26,8'h16,8'h24,8'h8d,8'h88,8'h64,8'h88,8'h72,8'h1c,8'h1b,8'h29,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h27,8'h25,8'h00,8'h3c,8'h98,8'h5a,8'h25,8'h41,8'h57,8'h63,8'h69,8'h6d,8'h73,8'h79,8'h76,8'h77,8'h76,8'h70,8'h6e,8'h6e,8'h67,8'h62,8'h54,8'h41,8'h33,8'h42,8'h6f,8'h9b,8'h8c,8'h58,8'h0d,8'h0b,8'h66,8'h31,8'h45,8'h68,8'h6a,8'h67,8'h53,8'h3e,8'h35,8'h53,8'h93,8'haa,8'h76,8'h3a,8'h00,8'h0b,8'h25,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h25,8'h0b,8'h6c,8'ha4,8'h80,8'h67,8'h66,8'h75,8'h8b,8'h8f,8'h7b,8'h54,8'h28,8'h02,8'h20,8'h25,8'h27,8'h23,8'h25,8'h8e,8'hb2,8'h9f,8'h4f,8'h1d,8'h24,8'h26,8'h27,8'h00,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h03,8'h55,8'h73,8'h32,8'h4f,8'h90,8'haf,8'h76,8'h2e,8'h17,8'h24,8'h27,8'h27,8'h00,8'h00,8'h27,8'h27,8'h22,8'h2e,8'h7c,8'h93,8'h89,8'h8b,8'h89,8'h73,8'h5f,8'h3f,8'h22,8'h11,8'h22,8'h27,8'h28,8'h27,8'h27,8'h11,8'h65,8'h81,8'h8a,8'h69,8'h1e,8'h21,8'h29,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h0c,8'h00,8'h00,8'h1d,8'h24,8'h25,8'h26,8'h26,8'h26,8'h25,8'h0c,8'h00,8'h38,8'h76,8'h98,8'h96,8'h2c,8'h00,8'h37,8'h75,8'h3c,8'h3f,8'h6b,8'h81,8'h89,8'h8c,8'h8c,8'h88,8'h88,8'h82,8'h79,8'h66,8'h3a,8'h47,8'ha1,8'h47,8'h00,8'h00,8'h45,8'h6b,8'h73,8'h75,8'h72,8'h5f,8'h44,8'h23,8'h00,8'h07,8'h23,8'h29,8'h27,8'h26,8'h23,8'h00,8'h45,8'h8a,8'h98,8'h69,8'h22,8'h0d,8'h29,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h27,8'h26,8'h0c,8'h00,8'h68,8'h98,8'h4b,8'h25,8'h33,8'h4a,8'h55,8'h63,8'h68,8'h6a,8'h6b,8'h69,8'h68,8'h64,8'h61,8'h5a,8'h4d,8'h3f,8'h38,8'h46,8'h6f,8'h99,8'h95,8'h69,8'h28,8'h00,8'h00,8'h3b,8'h69,8'h2b,8'h4e,8'h63,8'h57,8'h42,8'h33,8'h4f,8'h80,8'h99,8'h7e,8'h40,8'h00,8'h08,8'h23,8'h26,8'h00,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h11,8'h09,8'h45,8'h61,8'h69,8'h65,8'h53,8'h45,8'h2e,8'h20,8'h20,8'h23,8'h26,8'h27,8'h27,8'h00,8'h25,8'h03,8'h3a,8'h53,8'h38,8'h20,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h27,8'h27,8'h22,8'h2b,8'h83,8'h9d,8'haa,8'h89,8'h48,8'h1d,8'h25,8'h28,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h20,8'h21,8'h3d,8'h39,8'h2b,8'h23,8'h20,8'h1f,8'h21,8'h25,8'h27,8'h27,8'h00,8'h27,8'h27,8'h27,8'h20,8'h2f,8'h6b,8'h59,8'h23,8'h23,8'h28,8'h27,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h0d,8'h22,8'h27,8'h26,8'h27,8'h00,8'h27,8'h27,8'h26,8'h1b,8'h00,8'h31,8'h6d,8'h4e,8'h8a,8'h6a,8'h00,8'h00,8'h00,8'h52,8'h5c,8'h2b,8'h5f,8'h7d,8'h85,8'h8a,8'h8a,8'h88,8'h85,8'h83,8'h7a,8'h6b,8'h49,8'h32,8'h96,8'h57,8'h00,8'h00,8'h00,8'h0f,8'h24,8'h1d,8'h00,8'h00,8'h00,8'h19,8'h24,8'h28,8'h28,8'h00,8'h27,8'h00,8'h26,8'h23,8'h00,8'h0a,8'h20,8'h04,8'h20,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h22,8'h00,8'h1f,8'h73,8'h9e,8'h65,8'h2d,8'h25,8'h2e,8'h3a,8'h44,8'h4b,8'h50,8'h4d,8'h4a,8'h43,8'h39,8'h32,8'h43,8'h5d,8'h82,8'ha8,8'ha3,8'h76,8'h3b,8'h00,8'h00,8'h00,8'h00,8'h55,8'h4c,8'h29,8'h47,8'h40,8'h32,8'h4b,8'h89,8'ha8,8'h76,8'h3d,8'h00,8'h05,8'h24,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h24,8'h11,8'h10,8'h17,8'h10,8'h09,8'h0e,8'h23,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h25,8'h1f,8'h1f,8'h24,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h27,8'h27,8'h1b,8'h3c,8'h60,8'h4f,8'h26,8'h18,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h28,8'h26,8'h26,8'h24,8'h24,8'h25,8'h27,8'h27,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h23,8'h00,8'h00,8'h09,8'h25,8'h28,8'h27,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h28,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h21,8'h00,8'h22,8'h71,8'h47,8'h51,8'h93,8'h36,8'h00,8'h16,8'h00,8'h22,8'h6d,8'h32,8'h47,8'h77,8'h84,8'h89,8'h89,8'h8a,8'h88,8'h84,8'h7d,8'h70,8'h52,8'h33,8'h95,8'h5b,8'h00,8'h1d,8'h26,8'h24,8'h20,8'h1e,8'h1a,8'h23,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h25,8'h22,8'h21,8'h26,8'h28,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h26,8'h24,8'h00,8'h0f,8'h64,8'h8f,8'h84,8'h6a,8'h46,8'h38,8'h3e,8'h43,8'h44,8'h41,8'h3f,8'h44,8'h5b,8'h7d,8'h9e,8'ha9,8'h9b,8'h72,8'h3b,8'h00,8'h00,8'h0c,8'h20,8'h00,8'h00,8'h6b,8'h30,8'h25,8'h3c,8'h46,8'h75,8'h97,8'h8a,8'h4c,8'h0f,8'h0b,8'h22,8'h25,8'h28,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h28,8'h27,8'h27,8'h2a,8'h29,8'h28,8'h26,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h27,8'h28,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h27,8'h28,8'h20,8'h01,8'h0a,8'h24,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h28,8'h27,8'h00,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h24,8'h26,8'h26,8'h26,8'h27,8'h00,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h22,8'h00,8'h1a,8'h64,8'h4d,8'h2a,8'h83,8'h6e,8'h00,8'h13,8'h27,8'h20,8'h00,8'h69,8'h50,8'h35,8'h6c,8'h80,8'h88,8'h8b,8'h8c,8'h8a,8'h82,8'h7e,8'h74,8'h57,8'h35,8'h93,8'h57,8'h00,8'h1b,8'h27,8'h27,8'h28,8'h28,8'h27,8'h26,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h28,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h25,8'h1e,8'h00,8'h1d,8'h44,8'h71,8'h89,8'h97,8'ha0,8'ha4,8'ha3,8'ha3,8'ha0,8'h9c,8'h94,8'h82,8'h62,8'h3c,8'h21,8'h00,8'h00,8'h1d,8'h26,8'h26,8'h26,8'h09,8'h3a,8'h71,8'h38,8'h65,8'h98,8'h8d,8'h65,8'h36,8'h23,8'h17,8'h24,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h26,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h21,8'h00,8'h1f,8'h6e,8'h4f,8'h20,8'h57,8'h96,8'h33,8'h00,8'h25,8'h27,8'h24,8'h00,8'h55,8'h6d,8'h2c,8'h60,8'h81,8'h89,8'h8b,8'h8a,8'h8a,8'h85,8'h7e,8'h73,8'h4f,8'h36,8'h97,8'h48,8'h00,8'h24,8'h00,8'h27,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h22,8'h00,8'h00,8'h00,8'h21,8'h37,8'h4f,8'h60,8'h63,8'h5c,8'h4c,8'h3c,8'h25,8'h00,8'h00,8'h00,8'h12,8'h23,8'h26,8'h27,8'h27,8'h27,8'h25,8'h00,8'h61,8'ha9,8'ha3,8'ha2,8'h6a,8'h2e,8'h00,8'h1e,8'h27,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h21,8'h00,8'h0c,8'h6f,8'h60,8'h22,8'h29,8'h89,8'h6d,8'h00,8'h12,8'h26,8'h27,8'h22,8'h00,8'h52,8'h77,8'h2f,8'h5e,8'h7c,8'h87,8'h88,8'h89,8'h88,8'h81,8'h7c,8'h6e,8'h43,8'h4a,8'ha0,8'h30,8'h00,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h24,8'h20,8'h17,8'h0d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0a,8'h0b,8'h1b,8'h22,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h24,8'h0c,8'h6a,8'h93,8'h6b,8'h38,8'h0e,8'h1f,8'h26,8'h29,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h23,8'h00,8'h28,8'h67,8'h60,8'h2b,8'h22,8'h5f,8'h93,8'h2e,8'h00,8'h24,8'h26,8'h20,8'h0b,8'h38,8'h6d,8'h4f,8'h34,8'h68,8'h7d,8'h82,8'h84,8'h84,8'h81,8'h7d,8'h75,8'h63,8'h31,8'h67,8'h89,8'h0d,8'h22,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h26,8'h27,8'h25,8'h26,8'h24,8'h25,8'h27,8'h26,8'h27,8'h26,8'h26,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h26,8'h22,8'h00,8'h27,8'h21,8'h00,8'h19,8'h26,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h22,8'h00,8'h2c,8'h75,8'h55,8'h2c,8'h2e,8'h37,8'h91,8'h5f,8'h00,8'h13,8'h25,8'h08,8'h00,8'h50,8'h7b,8'h4a,8'h2e,8'h55,8'h75,8'h84,8'h86,8'h88,8'h87,8'h81,8'h7d,8'h71,8'h4f,8'h2d,8'h8d,8'h5c,8'h00,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h27,8'h27,8'h00,8'h27,8'h00,8'h27,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h10,8'h00,8'h00,8'h1c,8'h26,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h24,8'h00,8'h29,8'h75,8'h5b,8'h2b,8'h41,8'h31,8'h63,8'h87,8'h19,8'h00,8'h00,8'h02,8'h0f,8'h65,8'h7b,8'h44,8'h31,8'h54,8'h72,8'h7d,8'h85,8'h89,8'h88,8'h86,8'h7d,8'h75,8'h66,8'h39,8'h50,8'h8e,8'h29,8'h18,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h20,8'h27,8'h26,8'h26,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h22,8'h03,8'h45,8'h75,8'h56,8'h37,8'h46,8'h39,8'h41,8'h88,8'h4a,8'h00,8'h00,8'h00,8'h48,8'h67,8'h59,8'h3e,8'h41,8'h5c,8'h71,8'h7c,8'h84,8'h84,8'h83,8'h81,8'h7f,8'h75,8'h67,8'h45,8'h38,8'h84,8'h54,8'h00,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h20,8'h00,8'h4a,8'h81,8'h49,8'h2e,8'h4a,8'h48,8'h2a,8'h70,8'h6d,8'h00,8'h00,8'h22,8'h68,8'h78,8'h42,8'h2b,8'h48,8'h62,8'h71,8'h7a,8'h7c,8'h80,8'h81,8'h7e,8'h7b,8'h73,8'h68,8'h4d,8'h2b,8'h6a,8'h7a,8'h04,8'h21,8'h28,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h1a,8'h09,8'h4e,8'h80,8'h4c,8'h32,8'h4b,8'h51,8'h36,8'h4a,8'h88,8'h3d,8'h00,8'h47,8'h70,8'h67,8'h3c,8'h33,8'h51,8'h67,8'h72,8'h79,8'h80,8'h7e,8'h7d,8'h7e,8'h7b,8'h71,8'h66,8'h53,8'h32,8'h4f,8'h86,8'h39,8'h00,8'h25,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h16,8'h29,8'h71,8'h69,8'h3c,8'h3e,8'h54,8'h5a,8'h3f,8'h37,8'h86,8'h66,8'h53,8'h73,8'h5d,8'h3b,8'h39,8'h49,8'h5c,8'h6a,8'h72,8'h74,8'h7c,8'h80,8'h7a,8'h7a,8'h78,8'h72,8'h66,8'h4a,8'h30,8'h64,8'h84,8'h41,8'h00,8'h24,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h25,8'h00,8'h2e,8'h81,8'h73,8'h2d,8'h37,8'h54,8'h62,8'h53,8'h2d,8'h67,8'ha5,8'h8b,8'h76,8'h47,8'h29,8'h3c,8'h5a,8'h69,8'h6c,8'h72,8'h77,8'h7a,8'h7b,8'h7e,8'h79,8'h78,8'h6d,8'h62,8'h47,8'h2b,8'h60,8'h8e,8'h40,8'h00,8'h24,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h03,8'h33,8'h75,8'h69,8'h31,8'h38,8'h55,8'h61,8'h65,8'h41,8'h3f,8'h84,8'h80,8'h5d,8'h38,8'h33,8'h4a,8'h63,8'h6e,8'h75,8'h77,8'h78,8'h7a,8'h7c,8'h7b,8'h77,8'h72,8'h6e,8'h5c,8'h43,8'h3d,8'h62,8'h81,8'h41,8'h00,8'h21,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h25,8'h00,8'h61,8'h65,8'h2b,8'h42,8'h57,8'h66,8'h6b,8'h69,8'h34,8'h29,8'h3e,8'h32,8'h3f,8'h53,8'h64,8'h6b,8'h73,8'h79,8'h7a,8'h7a,8'h7d,8'h7c,8'h78,8'h76,8'h6d,8'h65,8'h56,8'h36,8'h3a,8'h81,8'h73,8'h2a,8'h00,8'h23,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h25,8'h00,8'h59,8'h52,8'h2d,8'h53,8'h61,8'h6a,8'h75,8'h73,8'h4a,8'h2b,8'h3d,8'h55,8'h66,8'h70,8'h74,8'h79,8'h7e,8'h7e,8'h7e,8'h7e,8'h81,8'h7d,8'h74,8'h6e,8'h66,8'h56,8'h3a,8'h40,8'h83,8'h73,8'h20,8'h00,8'h23,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h25,8'h00,8'h53,8'h59,8'h2c,8'h53,8'h63,8'h6d,8'h77,8'h79,8'h73,8'h6d,8'h6d,8'h71,8'h77,8'h7c,8'h7e,8'h7d,8'h7e,8'h7e,8'h7e,8'h7b,8'h77,8'h70,8'h6a,8'h61,8'h4c,8'h3c,8'h5a,8'h80,8'h63,8'h13,8'h05,8'h24,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h25,8'h00,8'h45,8'h5f,8'h2f,8'h53,8'h62,8'h6c,8'h76,8'h7c,8'h78,8'h7a,8'h79,8'h77,8'h7b,8'h7c,8'h7b,8'h7b,8'h7c,8'h7c,8'h79,8'h71,8'h6b,8'h64,8'h59,8'h42,8'h31,8'h6a,8'h8b,8'h44,8'h00,8'h12,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h25,8'h00,8'h39,8'h65,8'h32,8'h4e,8'h61,8'h6d,8'h76,8'h79,8'h7b,8'h7e,8'h7d,8'h7f,8'h7f,8'h7b,8'h79,8'h7a,8'h7b,8'h77,8'h71,8'h69,8'h63,8'h54,8'h40,8'h34,8'h6a,8'h85,8'h3b,8'h00,8'h12,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h00,8'h2a,8'h66,8'h30,8'h4a,8'h61,8'h6b,8'h75,8'h79,8'h7c,8'h7e,8'h7c,8'h7e,8'h7e,8'h7a,8'h77,8'h73,8'h73,8'h6d,8'h65,8'h60,8'h4c,8'h32,8'h50,8'h80,8'h63,8'h28,8'h00,8'h1b,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h00,8'h21,8'h65,8'h2e,8'h49,8'h5f,8'h68,8'h72,8'h77,8'h78,8'h78,8'h79,8'h7b,8'h7c,8'h76,8'h72,8'h6e,8'h6a,8'h64,8'h56,8'h44,8'h2e,8'h5b,8'h8e,8'h53,8'h00,8'h00,8'h24,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h26,8'h00,8'h21,8'h69,8'h30,8'h46,8'h59,8'h67,8'h6e,8'h75,8'h75,8'h79,8'h7b,8'h77,8'h77,8'h70,8'h6e,8'h65,8'h5d,8'h53,8'h3b,8'h37,8'h6c,8'h87,8'h45,8'h00,8'h03,8'h25,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h00,8'h19,8'h6a,8'h37,8'h43,8'h59,8'h65,8'h6d,8'h73,8'h73,8'h76,8'h76,8'h73,8'h6e,8'h69,8'h66,8'h5d,8'h4a,8'h33,8'h45,8'h7c,8'h79,8'h34,8'h00,8'h18,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h11,8'h02,8'h66,8'h3e,8'h41,8'h58,8'h65,8'h6a,8'h71,8'h72,8'h71,8'h6f,8'h6a,8'h67,8'h61,8'h53,8'h43,8'h2a,8'h51,8'h8f,8'h69,8'h19,8'h00,8'h21,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h1d,8'h00,8'h62,8'h40,8'h3f,8'h58,8'h62,8'h67,8'h6e,8'h6e,8'h6c,8'h66,8'h61,8'h58,8'h46,8'h38,8'h37,8'h5f,8'h88,8'h55,8'h05,8'h00,8'h25,8'h28,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1d,8'h00,8'h63,8'h41,8'h38,8'h54,8'h60,8'h66,8'h69,8'h65,8'h61,8'h58,8'h4c,8'h35,8'h2f,8'h5a,8'h7a,8'h5e,8'h2a,8'h00,8'h25,8'h28,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1c,8'h00,8'h63,8'h40,8'h35,8'h50,8'h59,8'h61,8'h61,8'h5b,8'h50,8'h46,8'h2e,8'h34,8'h70,8'h81,8'h46,8'h00,8'h00,8'h23,8'h28,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1f,8'h00,8'h63,8'h3f,8'h32,8'h4c,8'h54,8'h59,8'h55,8'h49,8'h37,8'h34,8'h4a,8'h7a,8'h6e,8'h29,8'h00,8'h10,8'h25,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h00,8'h64,8'h41,8'h33,8'h47,8'h4d,8'h4d,8'h3d,8'h28,8'h42,8'h7c,8'h74,8'h33,8'h00,8'h00,8'h25,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h19,8'h00,8'h63,8'h41,8'h2d,8'h42,8'h43,8'h32,8'h2f,8'h5b,8'h86,8'h5f,8'h0b,8'h00,8'h12,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1c,8'h00,8'h65,8'h3e,8'h26,8'h29,8'h2e,8'h53,8'h6a,8'h67,8'h40,8'h00,8'h00,8'h1e,8'h26,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1c,8'h0a,8'h68,8'h37,8'h18,8'h37,8'h70,8'h74,8'h33,8'h00,8'h00,8'h21,8'h29,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h1b,8'h72,8'h4d,8'h48,8'h7f,8'h5e,8'h1c,8'h00,8'h09,8'h24,8'h27,8'h00,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h1d,8'h88,8'h85,8'h55,8'h31,8'h00,8'h0a,8'h25,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h21,8'h06,8'h4e,8'h3e,8'h00,8'h00,8'h20,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h18,8'h00,8'h00,8'h00,8'h07,8'h24,8'h27,8'h00,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h0e,8'h00,8'h16,8'h27,8'h28,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h21,8'h27,8'h29,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h2a,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}};

parameter bit [7:0] SpriteTableB[111:0][226:0] = '{'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h27,8'h26,8'h26,8'h27,8'h27,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h26,8'h26,8'h25,8'h25,8'h21,8'h20,8'h1f,8'h1c,8'h15,8'h11,8'h11,8'h12,8'h0b,8'h08,8'h0a,8'h0b,8'h0e,8'h0d,8'h0b,8'h0b,8'h0b,8'h0c,8'h0c,8'h0b,8'h0a,8'h0e,8'h18,8'h20,8'h20,8'h1f,8'h1f,8'h24,8'h27,8'h25,8'h26,8'h26,8'h26,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h25,8'h22,8'h22,8'h23,8'h22,8'h11,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h02,8'h1e,8'h22,8'h22,8'h23,8'h23,8'h24,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h00,8'h26,8'h24,8'h23,8'h22,8'h1a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h12,8'h20,8'h23,8'h25,8'h26,8'h26,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h25,8'h24,8'h20,8'h12,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h08,8'h04,8'h04,8'h1f,8'h1f,8'h1b,8'h23,8'h24,8'h23,8'h25,8'h26,8'h28,8'h28,8'h27,8'h2a,8'h2a,8'h2b,8'h2c,8'h27,8'h26,8'h27,8'h26,8'h26,8'h26,8'h24,8'h21,8'h20,8'h22,8'h20,8'h10,8'h0a,8'h07,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0b,8'h1f,8'h22,8'h24,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h24,8'h20,8'h1a,8'h05,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'h10,8'h1f,8'h24,8'h22,8'h27,8'h2c,8'h31,8'h37,8'h41,8'h45,8'h43,8'h46,8'h4b,8'h4e,8'h4f,8'h4f,8'h4e,8'h4f,8'h51,8'h54,8'h50,8'h50,8'h50,8'h4f,8'h4e,8'h50,8'h51,8'h4e,8'h4d,8'h4b,8'h4d,8'h4c,8'h47,8'h41,8'h3c,8'h3c,8'h37,8'h2a,8'h27,8'h23,8'h1e,8'h0d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h13,8'h22,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h00,8'h26,8'h25,8'h23,8'h1a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0c,8'h16,8'h18,8'h23,8'h2c,8'h33,8'h3d,8'h43,8'h45,8'h45,8'h49,8'h4d,8'h4c,8'h4e,8'h4a,8'h4c,8'h4b,8'h4b,8'h4c,8'h4c,8'h4d,8'h49,8'h49,8'h49,8'h4a,8'h4c,8'h49,8'h43,8'h44,8'h45,8'h45,8'h44,8'h49,8'h49,8'h49,8'h4a,8'h4e,8'h4e,8'h4e,8'h50,8'h56,8'h59,8'h52,8'h4d,8'h50,8'h4c,8'h47,8'h42,8'h35,8'h28,8'h20,8'h17,8'h0e,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h1a,8'h22,8'h25,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h26,8'h25,8'h22,8'h10,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h05,8'h16,8'h24,8'h2c,8'h35,8'h40,8'h43,8'h46,8'h4b,8'h4a,8'h4a,8'h4a,8'h4d,8'h4c,8'h4d,8'h47,8'h45,8'h41,8'h3a,8'h33,8'h2e,8'h2c,8'h29,8'h26,8'h25,8'h24,8'h21,8'h1c,8'h1b,8'h1f,8'h1b,8'h1d,8'h1d,8'h1b,8'h18,8'h18,8'h1c,8'h19,8'h20,8'h23,8'h25,8'h27,8'h2c,8'h35,8'h3b,8'h3e,8'h41,8'h4a,8'h4f,8'h53,8'h56,8'h54,8'h52,8'h4e,8'h4d,8'h46,8'h40,8'h3c,8'h2a,8'h22,8'h0e,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1e,8'h23,8'h25,8'h26,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h25,8'h25,8'h22,8'h12,8'h06,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0b,8'h20,8'h26,8'h2d,8'h31,8'h36,8'h44,8'h4b,8'h4c,8'h51,8'h4e,8'h4b,8'h48,8'h43,8'h3d,8'h34,8'h34,8'h2f,8'h2b,8'h26,8'h1f,8'h13,8'h0c,8'h13,8'h06,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h00,8'h00,8'h00,8'h00,8'h12,8'h1e,8'h25,8'h2c,8'h34,8'h3f,8'h3a,8'h41,8'h49,8'h4a,8'h50,8'h4e,8'h4a,8'h44,8'h3c,8'h39,8'h2b,8'h1b,8'h10,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h26,8'h25,8'h25,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h23,8'h08,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h13,8'h23,8'h2e,8'h3f,8'h47,8'h4d,8'h4f,8'h52,8'h4f,8'h4d,8'h4b,8'h43,8'h40,8'h33,8'h29,8'h24,8'h1b,8'h0a,8'h02,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'h00,8'h05,8'h14,8'h1f,8'h25,8'h2d,8'h3b,8'h46,8'h4e,8'h59,8'h58,8'h4b,8'h45,8'h36,8'h28,8'h18,8'h03,8'h00,8'h00,8'h1b,8'h28,8'h00,8'h00,8'h21,8'h25,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h26,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h22,8'h0f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h09,8'h19,8'h23,8'h37,8'h42,8'h49,8'h53,8'h51,8'h4f,8'h4e,8'h4c,8'h4a,8'h44,8'h31,8'h27,8'h1e,8'h0f,8'h0c,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h09,8'h27,8'h21,8'h18,8'h21,8'h26,8'h24,8'h25,8'h1f,8'h2c,8'h27,8'h15,8'h13,8'h10,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h09,8'h19,8'h1e,8'h23,8'h2e,8'h3d,8'h4a,8'h55,8'h59,8'h53,8'h45,8'h2b,8'h1c,8'h1c,8'h20,8'h21,8'h00,8'h00,8'h00,8'h00,8'h20,8'h23,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h25,8'h24,8'h24,8'h21,8'h18,8'h19,8'h20,8'h24,8'h25,8'h26,8'h26,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h23,8'h1e,8'h02,8'h00,8'h00,8'h00,8'h00,8'h00,8'h17,8'h22,8'h33,8'h44,8'h4a,8'h4f,8'h55,8'h57,8'h54,8'h4d,8'h44,8'h35,8'h2b,8'h25,8'h1f,8'h05,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h18,8'h25,8'h2d,8'h3d,8'h43,8'h45,8'h45,8'h45,8'h46,8'h4a,8'h4e,8'h57,8'h51,8'h65,8'h61,8'h58,8'h56,8'h5d,8'h62,8'h68,8'h59,8'h68,8'h69,8'h5b,8'h5a,8'h56,8'h58,8'h4b,8'h53,8'h50,8'h40,8'h3e,8'h42,8'h43,8'h41,8'h38,8'h2f,8'h28,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h16,8'h24,8'h2a,8'h31,8'h42,8'h40,8'h2c,8'h3f,8'h53,8'h47,8'h34,8'h21,8'h00,8'h00,8'h00,8'h00,8'h00,8'h13,8'h23,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h00,8'h26,8'h24,8'h1f,8'h18,8'h0e,8'h03,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h05,8'h1f,8'h26,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h25,8'h21,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'h1d,8'h27,8'h3e,8'h4a,8'h56,8'h57,8'h53,8'h52,8'h49,8'h43,8'h31,8'h24,8'h17,8'h07,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h28,8'h31,8'h3e,8'h47,8'h4f,8'h51,8'h53,8'h55,8'h53,8'h53,8'h52,8'h51,8'h59,8'h69,8'h6b,8'h76,8'h62,8'h62,8'h63,8'h6f,8'h78,8'h51,8'h74,8'h87,8'h6e,8'h6c,8'h7f,8'h7c,8'h5e,8'h55,8'h55,8'h5f,8'h68,8'h6b,8'h58,8'h4c,8'h4e,8'h50,8'h51,8'h52,8'h56,8'h57,8'h54,8'h4f,8'h4b,8'h42,8'h2c,8'h1f,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h08,8'h2f,8'h48,8'h27,8'h36,8'h4d,8'h59,8'h58,8'h4b,8'h39,8'h24,8'h05,8'h00,8'h00,8'h00,8'h00,8'h10,8'h21,8'h25,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h22,8'h1d,8'h03,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h08,8'h00,8'h00,8'h00,8'h24,8'h26},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h25,8'h21,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h21,8'h25,8'h2f,8'h44,8'h51,8'h5a,8'h53,8'h4e,8'h46,8'h3d,8'h2e,8'h23,8'h14,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1b,8'h2a,8'h44,8'h4a,8'h47,8'h44,8'h39,8'h30,8'h2c,8'h3c,8'h45,8'h4f,8'h4d,8'h4d,8'h53,8'h55,8'h54,8'h54,8'h56,8'h5d,8'h6a,8'h71,8'h6e,8'h69,8'h64,8'h67,8'h67,8'h5d,8'h6a,8'h6f,8'h80,8'h76,8'h7d,8'h70,8'h57,8'h60,8'h65,8'h8c,8'hb7,8'hb7,8'h84,8'h62,8'h5c,8'h54,8'h58,8'h64,8'h62,8'h5d,8'h63,8'h6a,8'h67,8'h56,8'h51,8'h50,8'h4b,8'h4d,8'h46,8'h39,8'h23,8'h00,8'h00,8'h00,8'h00,8'h32,8'h5c,8'h35,8'h00,8'h0b,8'h20,8'h2d,8'h41,8'h51,8'h54,8'h4e,8'h45,8'h30,8'h24,8'h00,8'h00,8'h00,8'h00,8'h13,8'h24,8'h25,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h25,8'h24,8'h12,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0f,8'h1b,8'h22,8'h26,8'h23,8'h24,8'h24,8'h24,8'h26,8'h2a,8'h29,8'h24,8'h00,8'h00,8'h17,8'h26},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h22,8'h12,8'h00,8'h00,8'h00,8'h00,8'h00,8'h11,8'h27,8'h39,8'h47,8'h4e,8'h53,8'h58,8'h54,8'h4b,8'h3d,8'h29,8'h1f,8'h10,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1e,8'h2d,8'h3c,8'h4b,8'h71,8'h66,8'h5a,8'h5b,8'h47,8'h30,8'h00,8'h00,8'h00,8'h00,8'h00,8'h15,8'h47,8'h56,8'h51,8'h56,8'h58,8'h57,8'h55,8'h56,8'h5b,8'h60,8'h62,8'h6f,8'h63,8'h68,8'h63,8'h63,8'h64,8'h71,8'h5c,8'h60,8'h72,8'h7a,8'h68,8'h5a,8'h6c,8'h6d,8'h94,8'he7,8'hd3,8'h7e,8'h6d,8'h65,8'h58,8'h5a,8'h70,8'h7b,8'h63,8'h5a,8'h5d,8'h56,8'h55,8'h5b,8'h58,8'h55,8'h70,8'h81,8'h84,8'h67,8'h58,8'h4f,8'h31,8'h3c,8'h7a,8'h4c,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h21,8'h26,8'h33,8'h47,8'h52,8'h55,8'h4d,8'h33,8'h1b,8'h00,8'h00,8'h00,8'h00,8'h1a,8'h25,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h24,8'h1e,8'h00,8'h00,8'h00,8'h00,8'h0b,8'h17,8'h27,8'h30,8'h3d,8'h45,8'h4c,8'h52,8'h4d,8'h50,8'h54,8'h51,8'h53,8'h5b,8'h52,8'h26,8'h0c,8'h00,8'h00,8'h26},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h25,8'h15,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0d,8'h25,8'h40,8'h4e,8'h57,8'h5b,8'h57,8'h4d,8'h45,8'h30,8'h1f,8'h0a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h39,8'h4a,8'h4e,8'h4a,8'h4c,8'h4b,8'h53,8'h6b,8'h57,8'h41,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2c,8'h57,8'h4f,8'h55,8'h56,8'h56,8'h54,8'h55,8'h5b,8'h5c,8'h5c,8'h57,8'h55,8'h58,8'h5c,8'h59,8'h59,8'h63,8'h5d,8'h66,8'h63,8'h68,8'h61,8'h53,8'h59,8'h5c,8'h78,8'hae,8'ha7,8'h77,8'h57,8'h54,8'h54,8'h58,8'h5d,8'h69,8'h5e,8'h58,8'h53,8'h53,8'h74,8'h6d,8'h6e,8'h7a,8'h6a,8'h68,8'h6c,8'h5c,8'h79,8'h60,8'h44,8'h83,8'h68,8'h53,8'h45,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'h1e,8'h2c,8'h44,8'h57,8'h5c,8'h4c,8'h38,8'h21,8'h04,8'h00,8'h00,8'h00,8'h17,8'h24,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h23,8'h0b,8'h00,8'h00,8'h00,8'h07,8'h0a,8'h23,8'h2d,8'h44,8'h54,8'h53,8'h4d,8'h47,8'h3c,8'h36,8'h45,8'h5b,8'h66,8'h62,8'h66,8'h67,8'h5c,8'h27,8'h16,8'h00,8'h00,8'h26},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h26,8'h26,8'h26,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h24,8'h17,8'h00,8'h00,8'h00,8'h00,8'h03,8'h20,8'h2e,8'h3f,8'h4e,8'h5b,8'h5b,8'h56,8'h48,8'h41,8'h2e,8'h1f,8'h0d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1e,8'h2d,8'h53,8'h5f,8'h82,8'h76,8'h5a,8'h4f,8'h52,8'h52,8'h4b,8'h3e,8'h22,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h16,8'h4c,8'h51,8'h57,8'h5a,8'h57,8'h55,8'h58,8'h55,8'h54,8'h55,8'h55,8'h54,8'h56,8'h58,8'h58,8'h56,8'h56,8'h58,8'h5d,8'h58,8'h54,8'h58,8'h56,8'h59,8'h5a,8'h59,8'h75,8'h81,8'h71,8'h5c,8'h5b,8'h58,8'h57,8'h62,8'h68,8'h60,8'h58,8'h59,8'h5c,8'h7c,8'h6f,8'h7b,8'h84,8'h6c,8'h69,8'h6f,8'h66,8'h52,8'h55,8'h86,8'h70,8'h47,8'h69,8'h59,8'h57,8'h52,8'h3e,8'h2e,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h13,8'h1f,8'h31,8'h4c,8'h52,8'h4c,8'h3c,8'h2a,8'h06,8'h00,8'h00,8'h00,8'h0d,8'h21,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h25,8'h1f,8'h11,8'h00,8'h00,8'h00,8'h1a,8'h29,8'h30,8'h39,8'h47,8'h4b,8'h4a,8'h41,8'h2b,8'h1f,8'h16,8'h11,8'h12,8'h25,8'h50,8'h5f,8'h5a,8'h60,8'h62,8'h4b,8'h23,8'h00,8'h00,8'h02,8'h25},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h26,8'h25,8'h23,8'h23,8'h23,8'h21,8'h21,8'h24,8'h23,8'h26,8'h00,8'h26,8'h00,8'h00,8'h00,8'h00,8'h26,8'h25,8'h1a,8'h00,8'h00,8'h00,8'h00,8'h0a,8'h25,8'h3b,8'h4f,8'h5a,8'h56,8'h56,8'h54,8'h45,8'h2d,8'h1f,8'h0a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h3c,8'h44,8'h4a,8'h5a,8'h6b,8'h60,8'h51,8'h59,8'h52,8'h4b,8'h43,8'h2a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h17,8'h29,8'h2c,8'h0f,8'h00,8'h00,8'h00,8'h47,8'h56,8'h5f,8'h79,8'h6a,8'h63,8'h58,8'h51,8'h53,8'h55,8'h55,8'h55,8'h55,8'h55,8'h57,8'h55,8'h53,8'h54,8'h56,8'h56,8'h57,8'h59,8'h56,8'h59,8'h58,8'h4f,8'h68,8'h6f,8'h57,8'h5a,8'h6e,8'h5c,8'h54,8'h65,8'h67,8'h5b,8'h5a,8'h59,8'h5b,8'h61,8'h74,8'h71,8'h85,8'h6b,8'h75,8'h84,8'h44,8'h48,8'hae,8'h8d,8'h3b,8'h4d,8'h60,8'h59,8'h58,8'h59,8'h56,8'h57,8'h50,8'h48,8'h39,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0f,8'h23,8'h34,8'h4a,8'h51,8'h44,8'h28,8'h0f,8'h00,8'h00,8'h00,8'h0a,8'h24,8'h00,8'h00,8'h00,8'h26,8'h26,8'h24,8'h11,8'h00,8'h00,8'h0b,8'h22,8'h27,8'h3e,8'h55,8'h5e,8'h51,8'h3a,8'h25,8'h13,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h4c,8'h60,8'h5d,8'h63,8'h59,8'h2e,8'h1a,8'h00,8'h00,8'h23,8'h26},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h23,8'h1b,8'h0d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h17,8'h1f,8'h23,8'h26,8'h26,8'h25,8'h21,8'h00,8'h00,8'h00,8'h00,8'h05,8'h1d,8'h31,8'h4a,8'h57,8'h5a,8'h5c,8'h53,8'h45,8'h2d,8'h17,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'h33,8'h43,8'h4b,8'h4e,8'h4d,8'h53,8'h65,8'h62,8'h51,8'h4d,8'h51,8'h44,8'h2e,8'h03,8'h00,8'h00,8'h00,8'h00,8'h00,8'h08,8'h1f,8'h2a,8'h39,8'h47,8'h44,8'h1e,8'h00,8'h00,8'h00,8'h4e,8'h74,8'h7c,8'h79,8'h6d,8'h7b,8'h62,8'h59,8'h55,8'h54,8'h54,8'h54,8'h53,8'h54,8'h54,8'h55,8'h55,8'h56,8'h58,8'h58,8'h58,8'h57,8'h58,8'h59,8'h55,8'h58,8'h69,8'h61,8'h56,8'h59,8'h69,8'h5e,8'h55,8'h58,8'h59,8'h5a,8'h5b,8'h59,8'h5a,8'h65,8'h64,8'h5b,8'h6c,8'h69,8'h68,8'h52,8'h47,8'ha5,8'hab,8'h49,8'h48,8'h61,8'h65,8'h59,8'h5a,8'h5e,8'h5a,8'h55,8'h53,8'h79,8'h76,8'h56,8'h4c,8'h36,8'h02,8'h00,8'h00,8'h00,8'h00,8'h0c,8'h21,8'h31,8'h4a,8'h4c,8'h3f,8'h23,8'h01,8'h00,8'h00,8'h00,8'h1e,8'h25,8'h26,8'h25,8'h09,8'h00,8'h00,8'h00,8'h1a,8'h29,8'h3f,8'h51,8'h5a,8'h5d,8'h46,8'h26,8'h13,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h28,8'h56,8'h61,8'h66,8'h6f,8'h45,8'h18,8'h00,8'h00,8'h14,8'h27,8'h26},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h00,8'h23,8'h1f,8'h08,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'h28,8'h42,8'h4f,8'h59,8'h56,8'h54,8'h4b,8'h3b,8'h27,8'h13,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h14,8'h37,8'h42,8'h4e,8'h51,8'h51,8'h4f,8'h4f,8'h55,8'h54,8'h55,8'h52,8'h50,8'h47,8'h33,8'h1a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h13,8'h28,8'h37,8'h44,8'h48,8'h49,8'h4a,8'h47,8'h22,8'h00,8'h00,8'h00,8'h61,8'h67,8'h6c,8'h68,8'h6c,8'h99,8'h6a,8'h58,8'h58,8'h57,8'h55,8'h53,8'h52,8'h55,8'h5a,8'h59,8'h58,8'h57,8'h58,8'h57,8'h59,8'h59,8'h64,8'h72,8'h6b,8'h5d,8'h62,8'h5e,8'h65,8'h75,8'h6b,8'h5e,8'h58,8'h59,8'h5a,8'h5a,8'h59,8'h5a,8'h65,8'h6a,8'h62,8'h59,8'h5f,8'h5a,8'h46,8'h56,8'hb0,8'hac,8'h4a,8'h41,8'h52,8'h67,8'h73,8'h57,8'h50,8'h54,8'h54,8'h5c,8'h62,8'h6b,8'h63,8'h59,8'h61,8'h61,8'h66,8'h5a,8'h4a,8'h23,8'h00,8'h00,8'h00,8'h00,8'h1b,8'h2e,8'h3e,8'h44,8'h42,8'h2f,8'h07,8'h00,8'h00,8'h00,8'h05,8'h00,8'h00,8'h05,8'h1e,8'h2b,8'h43,8'h4d,8'h54,8'h59,8'h49,8'h2d,8'h13,8'h00,8'h00,8'h00,8'h00,8'h00,8'h09,8'h12,8'h00,8'h00,8'h0c,8'h33,8'h5d,8'h5d,8'h61,8'h55,8'h26,8'h00,8'h00,8'h00,8'h25,8'h26,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h0b,8'h14,8'h1a,8'h0d,8'h06,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h35,8'h4f,8'h5c,8'h5d,8'h5a,8'h52,8'h3b,8'h21,8'h0a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h18,8'h3b,8'h4c,8'h56,8'h59,8'h5b,8'h53,8'h51,8'h54,8'h51,8'h63,8'h5d,8'h52,8'h4b,8'h3e,8'h0d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h16,8'h27,8'h3d,8'h47,8'h47,8'h48,8'h49,8'h47,8'h49,8'h47,8'h21,8'h00,8'h00,8'h25,8'h73,8'h53,8'h58,8'h5f,8'h63,8'h6f,8'h5a,8'h54,8'h56,8'h54,8'h53,8'h52,8'h54,8'h59,8'h5f,8'h5f,8'h57,8'h54,8'h57,8'h55,8'h57,8'h68,8'h78,8'h7a,8'h76,8'h6a,8'h5e,8'h63,8'h63,8'h6e,8'h6a,8'h5c,8'h59,8'h59,8'h5a,8'h5b,8'h58,8'h59,8'h65,8'h6f,8'h63,8'h55,8'h52,8'h3e,8'h4e,8'hc2,8'hc7,8'h4a,8'h3a,8'h52,8'h5e,8'h72,8'h85,8'h59,8'h56,8'h53,8'h57,8'h5a,8'h59,8'h52,8'h5d,8'h7f,8'h82,8'h76,8'h90,8'h7e,8'h7a,8'h67,8'h49,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h23,8'h3e,8'h49,8'h3f,8'h29,8'h06,8'h00,8'h00,8'h00,8'h18,8'h27,8'h42,8'h56,8'h55,8'h55,8'h4f,8'h3d,8'h1f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1c,8'h23,8'h26,8'h26,8'h0c,8'h00,8'h1f,8'h4b,8'h5f,8'h5a,8'h57,8'h32,8'h11,8'h00,8'h00,8'h14,8'h26,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h21,8'h06,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h02,8'h16,8'h1c,8'h21,8'h2b,8'h35,8'h41,8'h49,8'h46,8'h44,8'h3c,8'h2a,8'h1f,8'h19,8'h07,8'h00,8'h00,8'h00,8'h20,8'h2e,8'h4e,8'h58,8'h58,8'h58,8'h53,8'h4b,8'h30,8'h0b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h39,8'h45,8'h4d,8'h50,8'h50,8'h55,8'h5a,8'h5f,8'h57,8'h59,8'h74,8'h65,8'h59,8'h4d,8'h44,8'h29,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0e,8'h1f,8'h32,8'h46,8'h4b,8'h49,8'h48,8'h48,8'h48,8'h48,8'h49,8'h45,8'h21,8'h00,8'h00,8'h20,8'h5a,8'h4d,8'h5a,8'h62,8'h57,8'h53,8'h55,8'h58,8'h56,8'h54,8'h59,8'h5a,8'h5a,8'h6d,8'h72,8'h69,8'h56,8'h56,8'h59,8'h5b,8'h5b,8'h65,8'h65,8'h62,8'h75,8'h71,8'h5f,8'h66,8'h59,8'h58,8'h59,8'h5a,8'h5a,8'h58,8'h5a,8'h5c,8'h5a,8'h59,8'h5f,8'h5e,8'h59,8'h51,8'h46,8'h56,8'hbe,8'hdd,8'h6b,8'h43,8'h57,8'h64,8'h7b,8'ha9,8'hb4,8'h85,8'h6a,8'h64,8'h6c,8'h6b,8'h55,8'h51,8'h63,8'h67,8'h6f,8'h88,8'h75,8'h78,8'h88,8'h78,8'h60,8'h65,8'h4c,8'h2f,8'h02,8'h00,8'h00,8'h00,8'h03,8'h21,8'h3e,8'h48,8'h32,8'h20,8'h1c,8'h24,8'h3c,8'h50,8'h53,8'h53,8'h53,8'h53,8'h42,8'h1d,8'h00,8'h00,8'h00,8'h00,8'h1e,8'h25,8'h26,8'h26,8'h26,8'h22,8'h00,8'h00,8'h28,8'h58,8'h5d,8'h5d,8'h43,8'h21,8'h00,8'h00,8'h00,8'h25,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h19,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h05,8'h1f,8'h2c,8'h42,8'h49,8'h4e,8'h4b,8'h51,8'h57,8'h5d,8'h59,8'h53,8'h56,8'h57,8'h4e,8'h4c,8'h49,8'h45,8'h30,8'h23,8'h31,8'h49,8'h4d,8'h55,8'h54,8'h51,8'h40,8'h29,8'h18,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h4c,8'h52,8'h69,8'h58,8'h52,8'h55,8'h70,8'h64,8'h5f,8'h57,8'h59,8'h5e,8'h60,8'h59,8'h47,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'h09,8'h0b,8'h20,8'h2e,8'h46,8'h47,8'h47,8'h48,8'h49,8'h48,8'h47,8'h45,8'h20,8'h00,8'h00,8'h05,8'h47,8'h51,8'h58,8'h59,8'h53,8'h50,8'h52,8'h55,8'h52,8'h5d,8'h70,8'h77,8'h6c,8'h6b,8'h69,8'h66,8'h5e,8'h66,8'h67,8'h64,8'h5f,8'h51,8'h55,8'h6a,8'h70,8'h5f,8'h55,8'h5c,8'h57,8'h56,8'h58,8'h5a,8'h5a,8'h5c,8'h5c,8'h5e,8'h60,8'h59,8'h65,8'h5f,8'h52,8'h43,8'h65,8'hce,8'he8,8'h78,8'h42,8'h61,8'h72,8'h89,8'hae,8'he8,8'hf1,8'hc0,8'h8a,8'h7e,8'h9f,8'h86,8'h63,8'h52,8'h54,8'h56,8'h5d,8'h72,8'h6d,8'h60,8'h6e,8'h6f,8'h59,8'h67,8'h67,8'h75,8'h63,8'h49,8'h2a,8'h00,8'h00,8'h00,8'h06,8'h25,8'h2d,8'h40,8'h48,8'h4c,8'h54,8'h56,8'h55,8'h52,8'h4b,8'h2d,8'h14,8'h00,8'h00,8'h00,8'h16,8'h24,8'h26,8'h26,8'h26,8'h26,8'h25,8'h00,8'h00,8'h22,8'h45,8'h63,8'h61,8'h48,8'h24,8'h00,8'h00,8'h00,8'h25,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h22,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h09,8'h20,8'h33,8'h44,8'h52,8'h5d,8'h5d,8'h5c,8'h52,8'h46,8'h3f,8'h36,8'h2e,8'h28,8'h27,8'h42,8'h55,8'h53,8'h53,8'h52,8'h54,8'h4c,8'h4d,8'h4d,8'h4e,8'h52,8'h49,8'h2b,8'h13,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2c,8'h4c,8'h6a,8'h5f,8'h57,8'h57,8'h54,8'h5a,8'h86,8'h6c,8'h60,8'h5c,8'h68,8'h65,8'h57,8'h46,8'h10,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h11,8'h3a,8'h4a,8'h47,8'h48,8'h48,8'h47,8'h46,8'h44,8'h21,8'h00,8'h00,8'h0f,8'h49,8'h52,8'h54,8'h55,8'h55,8'h53,8'h53,8'h52,8'h55,8'h66,8'h6d,8'h8a,8'h6b,8'h61,8'h64,8'h6f,8'h6a,8'h6c,8'h75,8'h68,8'h6a,8'h45,8'h32,8'h58,8'h5f,8'h54,8'h57,8'h59,8'h5a,8'h5b,8'h5d,8'h5a,8'h5b,8'h5f,8'h5f,8'h62,8'h70,8'h5f,8'h63,8'h5e,8'h41,8'h51,8'hc4,8'hfc,8'h9c,8'h3d,8'h4b,8'h5c,8'h5a,8'h5f,8'h84,8'hdd,8'he9,8'h9d,8'h62,8'h61,8'h6d,8'h67,8'h5e,8'h51,8'h53,8'h5e,8'h5f,8'h62,8'h75,8'h63,8'h5d,8'h6c,8'h60,8'h61,8'h63,8'h6b,8'h6b,8'h6a,8'h64,8'h51,8'h2b,8'h00,8'h00,8'h00,8'h00,8'h23,8'h40,8'h52,8'h55,8'h52,8'h50,8'h4b,8'h27,8'h0c,8'h00,8'h00,8'h00,8'h1b,8'h26,8'h26,8'h26,8'h26,8'h26,8'h26,8'h15,8'h00,8'h0d,8'h36,8'h57,8'h61,8'h50,8'h25,8'h01,8'h00,8'h00,8'h22,8'h26,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h19,8'h28,8'h37,8'h4a,8'h57,8'h5c,8'h57,8'h4c,8'h47,8'h36,8'h29,8'h22,8'h16,8'h03,8'h00,8'h06,8'h21,8'h44,8'h57,8'h52,8'h52,8'h54,8'h54,8'h4e,8'h4b,8'h4a,8'h49,8'h3d,8'h23,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h43,8'h52,8'h63,8'h56,8'h55,8'h58,8'h59,8'h59,8'h61,8'h65,8'h59,8'h6a,8'h6c,8'h71,8'h61,8'h64,8'h49,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0d,8'h2e,8'h46,8'h45,8'h47,8'h45,8'h45,8'h46,8'h45,8'h22,8'h00,8'h00,8'h0e,8'h48,8'h52,8'h57,8'h58,8'h5a,8'h5c,8'h5c,8'h5e,8'h64,8'h75,8'h72,8'h74,8'h5e,8'h62,8'h6b,8'h5b,8'h61,8'h67,8'h5c,8'h5f,8'h6a,8'h4d,8'h25,8'h3c,8'h53,8'h59,8'h56,8'h57,8'h5b,8'h5e,8'h5d,8'h5d,8'h5f,8'h60,8'h63,8'h63,8'h61,8'h66,8'h59,8'h49,8'h5c,8'hc0,8'hf7,8'hba,8'h4f,8'h47,8'h57,8'h5b,8'h5b,8'h58,8'h71,8'h99,8'hab,8'h7b,8'h5e,8'h54,8'h56,8'h58,8'h5e,8'h5e,8'h5c,8'h6f,8'h66,8'h6c,8'h81,8'h64,8'h5c,8'h66,8'h58,8'h5c,8'h67,8'h68,8'h69,8'h81,8'h7b,8'h80,8'h69,8'h41,8'h1a,8'h00,8'h00,8'h00,8'h0a,8'h29,8'h44,8'h4a,8'h4d,8'h2f,8'h09,8'h00,8'h00,8'h00,8'h16,8'h26,8'h26,8'h26,8'h26,8'h26,8'h26,8'h23,8'h00,8'h00,8'h29,8'h4c,8'h58,8'h4d,8'h2e,8'h12,8'h00,8'h00,8'h0f,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h23,8'h09,8'h00,8'h00,8'h00,8'h00,8'h17,8'h2b,8'h41,8'h59,8'h63,8'h60,8'h54,8'h47,8'h30,8'h1f,8'h11,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h29,8'h4e,8'h54,8'h50,8'h50,8'h55,8'h53,8'h50,8'h4d,8'h3a,8'h23,8'h0c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2f,8'h45,8'h4f,8'h59,8'h56,8'h56,8'h54,8'h55,8'h56,8'h59,8'h61,8'h67,8'h5d,8'h59,8'h6d,8'h6e,8'h77,8'h6b,8'h6c,8'h68,8'h50,8'h41,8'h54,8'h51,8'h3b,8'h36,8'h41,8'h41,8'h31,8'h20,8'h00,8'h00,8'h06,8'h2e,8'h49,8'h48,8'h46,8'h46,8'h45,8'h47,8'h44,8'h1f,8'h00,8'h00,8'h06,8'h50,8'h5e,8'h5c,8'h61,8'h6d,8'h6c,8'h6c,8'h77,8'h7c,8'h7d,8'h7d,8'h77,8'h59,8'h58,8'h5c,8'h5a,8'h5d,8'h61,8'h5e,8'h58,8'h56,8'h5c,8'h3b,8'h20,8'h43,8'h5b,8'h58,8'h5a,8'h5e,8'h55,8'h59,8'h63,8'h71,8'h71,8'h72,8'h72,8'h6b,8'h6a,8'h43,8'h64,8'hd2,8'hfa,8'hc0,8'h4d,8'h47,8'h5a,8'h5a,8'h5c,8'h5d,8'h59,8'h5c,8'h6c,8'h82,8'h58,8'h5b,8'h56,8'h56,8'h58,8'h5f,8'h67,8'h65,8'h80,8'h64,8'h5b,8'h62,8'h58,8'h58,8'h5c,8'h57,8'h5c,8'h6c,8'h61,8'h5f,8'h6c,8'h65,8'h62,8'h5d,8'h5a,8'h56,8'h4b,8'h30,8'h00,8'h00,8'h00,8'h0f,8'h24,8'h37,8'h33,8'h1f,8'h12,8'h27,8'h26,8'h27,8'h26,8'h26,8'h26,8'h26,8'h26,8'h25,8'h03,8'h00,8'h1e,8'h4b,8'h65,8'h5a,8'h2d,8'h13,8'h00,8'h00,8'h0a,8'h25,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h1e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h36,8'h54,8'h62,8'h63,8'h5b,8'h43,8'h28,8'h18,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h33,8'h51,8'h51,8'h4c,8'h4a,8'h4e,8'h4f,8'h44,8'h2e,8'h15,8'h1f,8'h22,8'h00,8'h00,8'h00,8'h0b,8'h41,8'h50,8'h59,8'h66,8'h69,8'h58,8'h54,8'h56,8'h58,8'h61,8'h62,8'h67,8'h5f,8'h5e,8'h63,8'h62,8'h5c,8'h6a,8'h67,8'h80,8'h85,8'h84,8'h66,8'h71,8'h75,8'h56,8'h5d,8'h6b,8'h6b,8'h62,8'h43,8'h00,8'h00,8'h07,8'h33,8'h4b,8'h47,8'h45,8'h47,8'h46,8'h48,8'h44,8'h1e,8'h00,8'h00,8'h24,8'h80,8'h75,8'h7f,8'h6a,8'h6e,8'h86,8'h7b,8'h6c,8'h6d,8'h6c,8'h7c,8'h6b,8'h54,8'h53,8'h57,8'h59,8'h59,8'h59,8'h5b,8'h5b,8'h56,8'h5e,8'h4a,8'h20,8'h26,8'h4c,8'h62,8'h63,8'h60,8'h41,8'h45,8'h6d,8'h86,8'h90,8'h81,8'h74,8'h61,8'h48,8'h5a,8'hc9,8'hfd,8'hde,8'h62,8'h3c,8'h52,8'h56,8'h5a,8'h5c,8'h59,8'h59,8'h5a,8'h6c,8'h7e,8'h5e,8'h62,8'h58,8'h5f,8'h61,8'h5c,8'h58,8'h56,8'h5b,8'h58,8'h58,8'h5a,8'h5b,8'h5b,8'h5a,8'h5a,8'h59,8'h5e,8'h5c,8'h59,8'h5d,8'h5b,8'h5c,8'h5b,8'h5d,8'h5c,8'h5f,8'h5c,8'h4b,8'h0b,8'h00,8'h00,8'h00,8'h1d,8'h2f,8'h3a,8'h26,8'h18,8'h24,8'h2c,8'h21,8'h24,8'h26,8'h26,8'h25,8'h07,8'h00,8'h0d,8'h38,8'h65,8'h63,8'h38,8'h10,8'h00,8'h00,8'h00,8'h24,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h00,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h47,8'h5d,8'h60,8'h5b,8'h4e,8'h2e,8'h1e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h10,8'h3e,8'h4f,8'h51,8'h4e,8'h4f,8'h4e,8'h46,8'h2a,8'h09,8'h00,8'h00,8'h00,8'h00,8'h00,8'h32,8'h4a,8'h53,8'h53,8'h5e,8'h6a,8'h64,8'h5a,8'h58,8'h58,8'h5f,8'h85,8'h66,8'h5f,8'h56,8'h59,8'h64,8'h56,8'h6e,8'h7f,8'h6c,8'h77,8'h74,8'h79,8'h66,8'h5b,8'h56,8'h6b,8'h78,8'h62,8'h64,8'h6e,8'h4e,8'h00,8'h00,8'h08,8'h35,8'h4c,8'h48,8'h47,8'h49,8'h48,8'h49,8'h48,8'h21,8'h00,8'h00,8'h29,8'h81,8'h70,8'h77,8'h6f,8'h64,8'h71,8'h76,8'h70,8'h77,8'h62,8'h64,8'h5e,8'h61,8'h62,8'h54,8'h57,8'h59,8'h59,8'h59,8'h5a,8'h59,8'h5c,8'h54,8'h38,8'h4c,8'h53,8'h8f,8'h85,8'h63,8'h30,8'h2b,8'h66,8'h6d,8'h6f,8'h6a,8'h5c,8'h3c,8'h50,8'hc0,8'hfd,8'hf1,8'h83,8'h3f,8'h50,8'h5a,8'h59,8'h59,8'h5b,8'h5b,8'h64,8'h75,8'h71,8'h84,8'h62,8'h61,8'h5e,8'h5e,8'h65,8'h80,8'h64,8'h55,8'h55,8'h57,8'h58,8'h5b,8'h5a,8'h5c,8'h5c,8'h5b,8'h5a,8'h59,8'h59,8'h5a,8'h5b,8'h5b,8'h5b,8'h5b,8'h5e,8'h63,8'h70,8'h73,8'h6c,8'h4e,8'h32,8'h00,8'h00,8'h00,8'h14,8'h29,8'h3c,8'h2d,8'h1e,8'h1f,8'h28,8'h26,8'h24,8'h26,8'h1f,8'h00,8'h00,8'h26,8'h58,8'h68,8'h45,8'h19,8'h00,8'h00,8'h00,8'h22,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h22,8'h00,8'h00,8'h00,8'h00,8'h15,8'h33,8'h53,8'h60,8'h5d,8'h51,8'h3f,8'h24,8'h06,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h34,8'h3f,8'h1f,8'h00,8'h00,8'h16,8'h42,8'h4d,8'h4d,8'h50,8'h4b,8'h39,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h10,8'h43,8'h5d,8'h64,8'h54,8'h52,8'h52,8'h55,8'h58,8'h57,8'h56,8'h59,8'h59,8'h5f,8'h62,8'h5b,8'h57,8'h52,8'h51,8'h5c,8'h81,8'h77,8'h6c,8'h75,8'h69,8'h68,8'h5e,8'h5c,8'h5e,8'h61,8'h73,8'h63,8'h67,8'h88,8'h51,8'h00,8'h00,8'h09,8'h32,8'h4b,8'h49,8'h4a,8'h4b,8'h48,8'h49,8'h47,8'h21,8'h00,8'h00,8'h3a,8'h78,8'h68,8'h64,8'h74,8'h6e,8'h6a,8'h6b,8'h8e,8'h76,8'h5a,8'h63,8'h6d,8'h81,8'h81,8'h59,8'h59,8'h5f,8'h5c,8'h59,8'h59,8'h5a,8'h5c,8'h61,8'h4a,8'h5d,8'h6d,8'h64,8'h75,8'h5f,8'h2e,8'h21,8'h52,8'h63,8'h5e,8'h60,8'h44,8'h4f,8'hbd,8'hf9,8'hf9,8'hab,8'h43,8'h4a,8'h58,8'h59,8'h5d,8'h5e,8'h5e,8'h5e,8'h61,8'h6b,8'h71,8'h80,8'h60,8'h5c,8'h5e,8'h59,8'h5b,8'h63,8'h5a,8'h57,8'h58,8'h60,8'h60,8'h59,8'h57,8'h5a,8'h59,8'h59,8'h59,8'h5c,8'h5b,8'h5a,8'h5c,8'h5e,8'h5e,8'h65,8'h6f,8'h69,8'h6a,8'h7f,8'h61,8'h59,8'h5a,8'h4c,8'h22,8'h00,8'h00,8'h01,8'h20,8'h38,8'h36,8'h22,8'h15,8'h27,8'h2d,8'h25,8'h00,8'h00,8'h1e,8'h45,8'h67,8'h4f,8'h23,8'h0e,8'h00,8'h00,8'h1f,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h23,8'h00,8'h00,8'h00,8'h00,8'h1f,8'h42,8'h59,8'h60,8'h63,8'h4f,8'h2e,8'h10,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h31,8'h48,8'h4d,8'h4d,8'h4d,8'h1f,8'h00,8'h00,8'h25,8'h4e,8'h51,8'h4d,8'h48,8'h2e,8'h13,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2c,8'h53,8'h6e,8'h5d,8'h5e,8'h57,8'h5d,8'h59,8'h55,8'h56,8'h59,8'h55,8'h5d,8'h5d,8'h54,8'h61,8'h5a,8'h53,8'h4d,8'h54,8'h61,8'h72,8'h69,8'h58,8'h73,8'h6d,8'h70,8'h69,8'h5e,8'h62,8'h5c,8'h7f,8'h66,8'h5e,8'h6c,8'h46,8'h00,8'h00,8'h07,8'h31,8'h4b,8'h4a,8'h4a,8'h4b,8'h4a,8'h4a,8'h44,8'h1f,8'h00,8'h00,8'h31,8'h70,8'h5f,8'h62,8'h63,8'h64,8'h59,8'h5a,8'h65,8'h5a,8'h5f,8'h5c,8'h6f,8'h7e,8'h6c,8'h54,8'h63,8'h7b,8'h75,8'h59,8'h5b,8'h5a,8'h5f,8'h6a,8'h64,8'h4c,8'h96,8'h58,8'h53,8'h5c,8'h3e,8'h3a,8'h4b,8'h5e,8'h5f,8'h4b,8'h47,8'hb2,8'hf8,8'hfd,8'hc6,8'h4e,8'h46,8'h59,8'h5b,8'h60,8'h62,8'h62,8'h61,8'h63,8'h5d,8'h67,8'h75,8'h70,8'h5d,8'h5a,8'h58,8'h58,8'h59,8'h56,8'h56,8'h66,8'h58,8'h68,8'h6a,8'h56,8'h56,8'h58,8'h59,8'h58,8'h59,8'h5f,8'h5e,8'h57,8'h5c,8'h60,8'h64,8'h66,8'h64,8'h72,8'h77,8'h6c,8'h66,8'h72,8'h65,8'h6f,8'h61,8'h3e,8'h00,8'h00,8'h00,8'h22,8'h29,8'h33,8'h24,8'h18,8'h29,8'h02,8'h00,8'h0d,8'h37,8'h5e,8'h53,8'h29,8'h19,8'h00,8'h00,8'h16,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h21,8'h00,8'h00,8'h00,8'h00,8'h28,8'h46,8'h5e,8'h60,8'h5c,8'h48,8'h28,8'h06,8'h00,8'h00,8'h00,8'h00,8'h21,8'h3c,8'h4a,8'h51,8'h51,8'h51,8'h54,8'h46,8'h00,8'h00,8'h00,8'h35,8'h53,8'h4d,8'h43,8'h2a,8'h11,8'h00,8'h00,8'h00,8'h00,8'h20,8'h3b,8'h51,8'h69,8'h79,8'h5f,8'h6d,8'h61,8'h58,8'h4f,8'h58,8'h66,8'h68,8'h55,8'h5e,8'h69,8'h74,8'h61,8'h57,8'h52,8'h65,8'h6d,8'h7e,8'h69,8'h5d,8'h59,8'h69,8'h6c,8'h80,8'h69,8'h5c,8'h5b,8'h59,8'h5c,8'h57,8'h54,8'h51,8'h42,8'h00,8'h00,8'h05,8'h35,8'h4a,8'h49,8'h48,8'h4a,8'h47,8'h4a,8'h47,8'h1f,8'h00,8'h00,8'h2e,8'h62,8'h55,8'h56,8'h56,8'h59,8'h56,8'h5e,8'h67,8'h59,8'h68,8'h6b,8'h6b,8'h6b,8'h63,8'h5e,8'h69,8'h73,8'h70,8'h59,8'h59,8'h5d,8'h63,8'h6f,8'h75,8'h4b,8'h77,8'ha5,8'h56,8'h46,8'h43,8'h65,8'h49,8'h51,8'h4b,8'h52,8'ha6,8'hf5,8'hfe,8'hd5,8'h63,8'h43,8'h5f,8'h63,8'h64,8'h65,8'h68,8'h61,8'h62,8'h63,8'h6d,8'h6d,8'h68,8'h5b,8'h58,8'h5b,8'h5e,8'h5b,8'h61,8'h64,8'h65,8'h7b,8'h5c,8'h59,8'h5d,8'h5e,8'h58,8'h55,8'h57,8'h58,8'h58,8'h5a,8'h63,8'h79,8'h68,8'h61,8'h63,8'h6d,8'h65,8'h6f,8'h81,8'h63,8'h60,8'h6d,8'h68,8'h78,8'h7d,8'h65,8'h46,8'h2c,8'h00,8'h00,8'h05,8'h23,8'h2b,8'h27,8'h20,8'h19,8'h1f,8'h2e,8'h54,8'h51,8'h2d,8'h11,8'h00,8'h00,8'h0a,8'h27,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h24,8'h00,8'h00,8'h00,8'h00,8'h2f,8'h55,8'h60,8'h5c,8'h5a,8'h43,8'h1f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h36,8'h4d,8'h55,8'h57,8'h55,8'h56,8'h58,8'h5c,8'h3d,8'h00,8'h00,8'h10,8'h41,8'h54,8'h3e,8'h1f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h34,8'h4b,8'h51,8'h53,8'h74,8'h7f,8'h5b,8'h76,8'h59,8'h33,8'h29,8'h52,8'h85,8'h6d,8'h51,8'h5a,8'h65,8'h85,8'h6b,8'h61,8'h5d,8'h8c,8'hc1,8'hd9,8'h97,8'h5e,8'h5d,8'h69,8'h63,8'h60,8'h5c,8'h5b,8'h59,8'h5a,8'h58,8'h58,8'h57,8'h55,8'h43,8'h00,8'h00,8'h03,8'h37,8'h4a,8'h4b,8'h4b,8'h51,8'h53,8'h4e,8'h49,8'h20,8'h00,8'h00,8'h1f,8'h4d,8'h56,8'h5c,8'h5b,8'h5e,8'h57,8'h5b,8'h64,8'h5b,8'h63,8'h80,8'h74,8'h71,8'h78,8'h78,8'h62,8'h58,8'h59,8'h5e,8'h5c,8'h61,8'h67,8'h77,8'h6a,8'h51,8'h46,8'hb6,8'ha5,8'h35,8'h2f,8'h83,8'h50,8'h38,8'h51,8'hbf,8'hf8,8'hfe,8'he1,8'h68,8'h3e,8'h58,8'h66,8'h6d,8'h6f,8'h69,8'h6a,8'h6a,8'h64,8'h5b,8'h68,8'h65,8'h5e,8'h5d,8'h68,8'h84,8'h6a,8'h5b,8'h66,8'h6d,8'h61,8'h66,8'h5a,8'h58,8'h58,8'h5a,8'h58,8'h57,8'h55,8'h53,8'h57,8'h58,8'h64,8'h82,8'h6a,8'h68,8'h60,8'h6d,8'h6c,8'h5e,8'h64,8'h67,8'h55,8'h54,8'h6a,8'h74,8'h72,8'h83,8'h66,8'h81,8'h54,8'h20,8'h00,8'h00,8'h08,8'h22,8'h28,8'h22,8'h2a,8'h4f,8'h55,8'h2c,8'h0b,8'h00,8'h00,8'h00,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h06,8'h00,8'h00,8'h0f,8'h2d,8'h57,8'h64,8'h60,8'h57,8'h42,8'h20,8'h00,8'h00,8'h00,8'h00,8'h26,8'h42,8'h4f,8'h51,8'h53,8'h55,8'h59,8'h68,8'h56,8'h51,8'h2d,8'h00,8'h00,8'h1d,8'h42,8'h38,8'h10,8'h00,8'h00,8'h00,8'h00,8'h07,8'h42,8'h4e,8'h51,8'h55,8'h58,8'h6c,8'h69,8'h4b,8'h36,8'h1a,8'h00,8'h31,8'h5a,8'h64,8'h63,8'h56,8'h5a,8'h60,8'h83,8'h6a,8'h64,8'h73,8'h98,8'he0,8'hf1,8'hb3,8'h72,8'h65,8'h69,8'h5e,8'h58,8'h58,8'h5a,8'h57,8'h57,8'h58,8'h5d,8'h5f,8'h63,8'h41,8'h00,8'h00,8'h06,8'h3c,8'h4b,8'h49,8'h4a,8'h4d,8'h4e,8'h4b,8'h45,8'h1f,8'h00,8'h00,8'h19,8'h4d,8'h58,8'h5a,8'h64,8'h63,8'h5a,8'h57,8'h59,8'h59,8'h67,8'h66,8'h79,8'h76,8'h61,8'h59,8'h59,8'h54,8'h63,8'h85,8'h71,8'h71,8'h7b,8'h8d,8'h67,8'h5b,8'h41,8'h7e,8'hdf,8'h7a,8'h38,8'ha0,8'h77,8'h43,8'hb4,8'hfb,8'hfe,8'hef,8'h89,8'h3d,8'h54,8'h68,8'h61,8'h5c,8'h52,8'h56,8'h71,8'h81,8'h65,8'h58,8'h60,8'h62,8'h62,8'h69,8'h6d,8'h90,8'h65,8'h5f,8'h61,8'h6a,8'h6a,8'h56,8'h54,8'h5a,8'h54,8'h55,8'h4f,8'h47,8'h36,8'h2b,8'h4d,8'h60,8'h63,8'h5e,8'h5c,8'h5d,8'h5a,8'h5b,8'h5a,8'h58,8'h5c,8'h61,8'h5e,8'h59,8'h6a,8'h80,8'h5f,8'h60,8'h62,8'h74,8'h62,8'h59,8'h37,8'h00,8'h00,8'h00,8'h21,8'h39,8'h4b,8'h53,8'h34,8'h14,8'h00,8'h00,8'h04,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h1e,8'h00,8'h00,8'h00,8'h1f,8'h39,8'h58,8'h66,8'h5a,8'h57,8'h42,8'h22,8'h00,8'h00,8'h00,8'h00,8'h33,8'h4d,8'h51,8'h55,8'h56,8'h58,8'h59,8'h6d,8'h76,8'h64,8'h53,8'h1b,8'h00,8'h00,8'h1f,8'h26,8'h09,8'h00,8'h00,8'h00,8'h00,8'h47,8'h57,8'h51,8'h51,8'h58,8'h55,8'h50,8'h46,8'h31,8'h00,8'h00,8'h00,8'h04,8'h56,8'h6c,8'h58,8'h59,8'h58,8'h59,8'h5b,8'h67,8'h61,8'h56,8'h5e,8'h76,8'h9b,8'hbd,8'h8a,8'h5a,8'h53,8'h56,8'h58,8'h57,8'h58,8'h5b,8'h58,8'h54,8'h5f,8'h68,8'h71,8'h73,8'h43,8'h00,8'h00,8'h0b,8'h3d,8'h4a,8'h4a,8'h46,8'h47,8'h45,8'h48,8'h46,8'h20,8'h00,8'h00,8'h28,8'h65,8'h61,8'h64,8'h67,8'h62,8'h5f,8'h64,8'h63,8'h5e,8'h5d,8'h5a,8'h69,8'h6c,8'h5c,8'h58,8'h5a,8'h5a,8'h66,8'h8a,8'h73,8'h6d,8'h6c,8'h6f,8'h63,8'h62,8'h4d,8'h46,8'hc2,8'hdc,8'h9a,8'hcf,8'hc8,8'hb7,8'hf3,8'hfd,8'hf4,8'h94,8'h37,8'h3e,8'h47,8'h43,8'h3e,8'h31,8'h2b,8'h4f,8'h71,8'h70,8'h62,8'h5c,8'h62,8'h67,8'h71,8'h63,8'h66,8'h6a,8'h5f,8'h79,8'h5d,8'h65,8'h63,8'h54,8'h51,8'h51,8'h46,8'h39,8'h28,8'h00,8'h00,8'h00,8'h5e,8'h66,8'h5e,8'h5b,8'h5a,8'h5b,8'h5b,8'h5b,8'h5c,8'h5f,8'h66,8'h75,8'h62,8'h5c,8'h5f,8'h66,8'h5d,8'h5e,8'h66,8'h79,8'h75,8'h75,8'h51,8'h00,8'h00,8'h00,8'h21,8'h48,8'h53,8'h35,8'h0f,8'h00,8'h00,8'h00,8'h24,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h22,8'h00,8'h00,8'h00,8'h1e,8'h32,8'h5b,8'h63,8'h61,8'h59,8'h46,8'h1d,8'h00,8'h00,8'h00,8'h00,8'h39,8'h4d,8'h54,8'h57,8'h58,8'h5a,8'h5a,8'h56,8'h63,8'h6a,8'h81,8'h4e,8'h00,8'h00,8'h09,8'h10,8'h00,8'h00,8'h00,8'h00,8'h00,8'h38,8'h5e,8'h58,8'h50,8'h53,8'h53,8'h38,8'h15,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3c,8'h57,8'h5b,8'h58,8'h58,8'h5a,8'h58,8'h58,8'h5b,8'h5e,8'h5b,8'h65,8'h6f,8'h6b,8'h80,8'h6b,8'h5d,8'h59,8'h59,8'h58,8'h54,8'h57,8'h5a,8'h57,8'h5f,8'h85,8'h85,8'h78,8'h76,8'h44,8'h00,8'h00,8'h0b,8'h40,8'h4d,8'h4b,8'h47,8'h4a,8'h47,8'h49,8'h46,8'h21,8'h00,8'h00,8'h26,8'h79,8'h7b,8'h6d,8'h5d,8'h5e,8'h61,8'h65,8'h60,8'h63,8'h5b,8'h5d,8'h5d,8'h58,8'h62,8'h6c,8'h6e,8'h68,8'h6a,8'h93,8'h85,8'h6a,8'h61,8'h5c,8'h62,8'h63,8'h5c,8'h33,8'h7b,8'hf2,8'hf9,8'hf9,8'hfb,8'hfe,8'hfd,8'hfd,8'hc4,8'h3c,8'h28,8'h46,8'h53,8'h41,8'h1e,8'h27,8'h46,8'h63,8'h62,8'h5c,8'h5f,8'h61,8'h6b,8'h6c,8'h73,8'h67,8'h64,8'h65,8'h5e,8'h6a,8'h5b,8'h58,8'h55,8'h52,8'h46,8'h30,8'h00,8'h00,8'h00,8'h00,8'h00,8'h39,8'h5e,8'h5a,8'h59,8'h58,8'h59,8'h5a,8'h5b,8'h60,8'h74,8'h6e,8'h6a,8'h86,8'h60,8'h5a,8'h5b,8'h5f,8'h63,8'h5e,8'h63,8'h6b,8'h76,8'h6d,8'h34,8'h00,8'h00,8'h1f,8'h39,8'h56,8'h36,8'h16,8'h00,8'h00,8'h00,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h25,8'h00,8'h00,8'h00,8'h1f,8'h36,8'h55,8'h62,8'h5d,8'h60,8'h55,8'h2a,8'h00,8'h00,8'h00,8'h00,8'h31,8'h52,8'h58,8'h58,8'h58,8'h58,8'h5e,8'h5c,8'h57,8'h58,8'h59,8'h65,8'h3b,8'h00,8'h00,8'h07,8'h00,8'h00,8'h00,8'h00,8'h07,8'h41,8'h51,8'h55,8'h48,8'h47,8'h40,8'h19,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1f,8'h53,8'h75,8'h5c,8'h57,8'h5b,8'h5c,8'h5a,8'h5b,8'h5d,8'h5d,8'h59,8'h5b,8'h5c,8'h67,8'h7d,8'h5a,8'h54,8'h5c,8'h5e,8'h5d,8'h60,8'h5b,8'h59,8'h5d,8'h69,8'h76,8'h72,8'h6c,8'h73,8'h41,8'h00,8'h00,8'h11,8'h46,8'h52,8'h4d,8'h4a,8'h4c,8'h49,8'h48,8'h44,8'h1f,8'h00,8'h00,8'h24,8'h65,8'h71,8'h64,8'h60,8'h75,8'h5c,8'h5b,8'h61,8'h6b,8'h6e,8'h67,8'h64,8'h5c,8'h6e,8'h85,8'h6a,8'h61,8'h61,8'h6c,8'h65,8'h55,8'h52,8'h4e,8'h4d,8'h48,8'h43,8'h30,8'h53,8'hde,8'hfd,8'hfd,8'hfd,8'hfb,8'hfb,8'hfb,8'hd4,8'h8e,8'h93,8'h8f,8'h59,8'h38,8'h41,8'h54,8'h62,8'h61,8'h5c,8'h5d,8'h5a,8'h61,8'h63,8'h69,8'h65,8'h62,8'h57,8'h5d,8'h61,8'h5f,8'h6b,8'h4b,8'h3f,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h4d,8'h57,8'h57,8'h57,8'h56,8'h59,8'h5c,8'h64,8'h69,8'h77,8'h6b,8'h62,8'h6f,8'h5f,8'h56,8'h60,8'h63,8'h6a,8'h68,8'h60,8'h5c,8'h5c,8'h47,8'h00,8'h00,8'h0d,8'h28,8'h4f,8'h40,8'h1e,8'h01,8'h00,8'h00,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h16,8'h00,8'h00,8'h13,8'h39,8'h5c,8'h63,8'h5c,8'h60,8'h5a,8'h34,8'h00,8'h00,8'h00,8'h00,8'h34,8'h50,8'h59,8'h59,8'h59,8'h59,8'h59,8'h68,8'h6c,8'h77,8'h6a,8'h60,8'h53,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h30,8'h53,8'h5c,8'h4c,8'h45,8'h28,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h45,8'h5d,8'h65,8'h58,8'h5a,8'h5c,8'h5d,8'h5a,8'h5b,8'h5e,8'h5e,8'h5b,8'h56,8'h51,8'h58,8'h68,8'h48,8'h49,8'h54,8'h65,8'h8a,8'h80,8'h75,8'h75,8'h7c,8'h83,8'h76,8'h67,8'h63,8'h6a,8'h41,8'h00,8'h00,8'h1a,8'h45,8'h4f,8'h4e,8'h4b,8'h4c,8'h49,8'h48,8'h44,8'h1e,8'h00,8'h00,8'h23,8'h51,8'h6c,8'h86,8'h83,8'h82,8'h6d,8'h6b,8'h91,8'h7c,8'h67,8'h69,8'h59,8'h37,8'h2d,8'h35,8'h28,8'h28,8'h2c,8'h43,8'h58,8'h65,8'h71,8'h7d,8'h81,8'h85,8'h92,8'ha0,8'hba,8'hf0,8'hfb,8'hfb,8'hfd,8'hfb,8'hfd,8'hfd,8'hf4,8'h99,8'h4c,8'h39,8'h30,8'h42,8'h52,8'h58,8'h5a,8'h57,8'h62,8'h72,8'h77,8'h7e,8'h5c,8'h5e,8'h5d,8'h5c,8'h55,8'h54,8'h43,8'h29,8'h29,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h21,8'h4c,8'h58,8'h56,8'h5d,8'h5b,8'h5d,8'h60,8'h64,8'h63,8'h69,8'h67,8'h5b,8'h72,8'h81,8'h6f,8'h57,8'h71,8'h6c,8'h6e,8'h70,8'h64,8'h5c,8'h44,8'h00,8'h00,8'h00,8'h25,8'h45,8'h34,8'h17,8'h00,8'h00,8'h00,8'h1f,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h17,8'h00,8'h00,8'h00,8'h2b,8'h5b,8'h66,8'h60,8'h5b,8'h5f,8'h44,8'h08,8'h00,8'h00,8'h00,8'h2b,8'h4d,8'h59,8'h58,8'h59,8'h5a,8'h5a,8'h5b,8'h5e,8'h6d,8'h80,8'h79,8'h63,8'h4b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h36,8'h6b,8'h54,8'h43,8'h23,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h37,8'h58,8'h6a,8'h6a,8'h55,8'h5d,8'h5d,8'h5d,8'h5f,8'h5e,8'h5a,8'h58,8'h4c,8'h32,8'h16,8'h00,8'h00,8'h00,8'h09,8'h2b,8'h43,8'h73,8'h81,8'h89,8'h85,8'h76,8'h6d,8'h65,8'h62,8'h68,8'h6d,8'h42,8'h00,8'h00,8'h1e,8'h45,8'h4e,8'h4c,8'h49,8'h48,8'h49,8'h4a,8'h44,8'h19,8'h00,8'h00,8'h24,8'h68,8'h5f,8'h76,8'h8b,8'h89,8'h78,8'h70,8'h6d,8'h69,8'h61,8'h5f,8'h61,8'h48,8'h3f,8'h2d,8'h20,8'h11,8'h15,8'h29,8'h42,8'h50,8'h65,8'h85,8'h94,8'ha6,8'hc7,8'hdb,8'hf6,8'hfb,8'hfa,8'hfb,8'hfd,8'hfb,8'hfd,8'hff,8'hf9,8'h9d,8'h4c,8'h43,8'h3f,8'h3d,8'h2f,8'h2a,8'h2c,8'h2b,8'h2f,8'h41,8'h5a,8'h67,8'h5a,8'h58,8'h50,8'h45,8'h30,8'h15,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h45,8'h58,8'h5b,8'h58,8'h5e,8'h5e,8'h63,8'h66,8'h6a,8'h7d,8'h6e,8'h68,8'h5d,8'h65,8'h76,8'h75,8'h64,8'h81,8'h83,8'h6f,8'h5f,8'h52,8'h46,8'h05,8'h00,8'h00,8'h20,8'h40,8'h40,8'h18,8'h00,8'h00,8'h00,8'h1a,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h21,8'h00,8'h00,8'h00,8'h27,8'h4c,8'h62,8'h62,8'h66,8'h61,8'h4f,8'h26,8'h00,8'h00,8'h00,8'h0f,8'h47,8'h58,8'h5b,8'h5b,8'h5a,8'h58,8'h59,8'h5d,8'h64,8'h70,8'h7c,8'h69,8'h58,8'h44,8'h00,8'h00,8'h00,8'h00,8'h00,8'h39,8'h4a,8'h43,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h29,8'h56,8'h62,8'h70,8'h70,8'h59,8'h5d,8'h5b,8'h56,8'h51,8'h46,8'h35,8'h21,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h47,8'h5e,8'h6a,8'h68,8'h56,8'h58,8'h5f,8'h7b,8'h85,8'h42,8'h00,8'h00,8'h1b,8'h46,8'h4d,8'h4a,8'h49,8'h4a,8'h4a,8'h4a,8'h43,8'h13,8'h00,8'h00,8'h2a,8'h81,8'h7d,8'h74,8'h80,8'h81,8'h6f,8'h74,8'h66,8'h62,8'h5c,8'h56,8'h57,8'h4c,8'h44,8'h2c,8'h00,8'h00,8'h00,8'h00,8'h05,8'h0a,8'h0e,8'h1f,8'h1f,8'h25,8'h44,8'h84,8'he8,8'hfd,8'hfb,8'hfd,8'hfd,8'hfb,8'he6,8'hbf,8'hb3,8'ha3,8'h8e,8'h82,8'h66,8'h4d,8'h35,8'h24,8'h22,8'h26,8'h28,8'h28,8'h39,8'h44,8'h42,8'h31,8'h19,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1f,8'h17,8'h0f,8'h00,8'h00,8'h00,8'h3e,8'h51,8'h58,8'h6a,8'h6a,8'h6a,8'h61,8'h63,8'h5e,8'h5c,8'h79,8'h79,8'h6a,8'h67,8'h6b,8'h63,8'h5d,8'h68,8'h62,8'h66,8'h5d,8'h35,8'h21,8'h00,8'h00,8'h00,8'h1f,8'h2f,8'h40,8'h23,8'h06,8'h00,8'h00,8'h00,8'h06,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h25,8'h00,8'h00,8'h00,8'h24,8'h4c,8'h65,8'h60,8'h5e,8'h61,8'h5f,8'h3d,8'h00,8'h00,8'h00,8'h00,8'h40,8'h57,8'h5a,8'h5c,8'h5d,8'h5d,8'h5b,8'h5d,8'h5d,8'h57,8'h5e,8'h6b,8'h59,8'h53,8'h32,8'h00,8'h00,8'h00,8'h00,8'h2e,8'h31,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h14,8'h23,8'h1a,8'h00,8'h00,8'h00,8'h00,8'h5e,8'h83,8'h76,8'h6c,8'h59,8'h52,8'h4e,8'h41,8'h21,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1a,8'h47,8'h5d,8'h58,8'h5a,8'h5f,8'h7d,8'h81,8'h3e,8'h00,8'h00,8'h14,8'h47,8'h4e,8'h48,8'h49,8'h4b,8'h48,8'h4b,8'h44,8'h11,8'h00,8'h00,8'h23,8'h69,8'h83,8'h79,8'h86,8'h80,8'h7c,8'h64,8'h5b,8'h4b,8'h3b,8'h23,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h06,8'h0a,8'h04,8'h09,8'h12,8'h2f,8'h57,8'h89,8'hdf,8'hfd,8'hfd,8'hfd,8'hfe,8'hfc,8'ha1,8'h3a,8'h3a,8'h43,8'h4a,8'h51,8'h5a,8'h56,8'h58,8'h58,8'h4b,8'h46,8'h3e,8'h28,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1a,8'h2e,8'h45,8'h30,8'h08,8'h00,8'h00,8'h00,8'h00,8'h41,8'h54,8'h5a,8'h66,8'h7d,8'h72,8'h5a,8'h5c,8'h5c,8'h68,8'h70,8'h8b,8'h6b,8'h79,8'h74,8'h4f,8'h4a,8'h42,8'h2b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0a,8'h2d,8'h34,8'h22,8'h17,8'h0e,8'h07,8'h00,8'h00,8'h00,8'h00,8'h23,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h18,8'h00,8'h00,8'h18,8'h3b,8'h62,8'h63,8'h63,8'h5e,8'h58,8'h53,8'h21,8'h00,8'h00,8'h00,8'h2c,8'h57,8'h5d,8'h5d,8'h5c,8'h5d,8'h5c,8'h5a,8'h5e,8'h71,8'h61,8'h5e,8'h5e,8'h52,8'h4c,8'h0a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h14,8'h27,8'h40,8'h34,8'h09,8'h00,8'h00,8'h00,8'h33,8'h5b,8'h79,8'h66,8'h4d,8'h41,8'h2e,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h09,8'h14,8'h12,8'h12,8'h13,8'h09,8'h00,8'h00,8'h00,8'h00,8'h00,8'h14,8'h4a,8'h5c,8'h5c,8'h5d,8'h5b,8'h60,8'h35,8'h00,8'h00,8'h18,8'h47,8'h4f,8'h49,8'h4a,8'h49,8'h47,8'h48,8'h45,8'h19,8'h00,8'h00,8'h27,8'h85,8'h7c,8'h76,8'h6b,8'h6f,8'h6f,8'h3b,8'h22,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h08,8'h1b,8'h24,8'h2a,8'h2b,8'h1f,8'h1f,8'h21,8'h29,8'h23,8'h30,8'hb4,8'hfe,8'hfb,8'hf9,8'hfa,8'hfc,8'ha3,8'h40,8'h4c,8'h5a,8'h6a,8'h69,8'h74,8'h82,8'h52,8'h3d,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1f,8'h28,8'h37,8'h48,8'h4f,8'h42,8'h1e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1b,8'h4e,8'h5b,8'h5a,8'h5f,8'h5c,8'h58,8'h57,8'h5b,8'h7c,8'h6a,8'h68,8'h5f,8'h52,8'h46,8'h31,8'h07,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h19,8'h25,8'h43,8'h2b,8'h29,8'h2d,8'h2f,8'h21,8'h0f,8'h01,8'h00,8'h00,8'h00,8'h24,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h21,8'h00,8'h00,8'h07,8'h2c,8'h54,8'h65,8'h62,8'h60,8'h5d,8'h56,8'h40,8'h00,8'h00,8'h00,8'h00,8'h49,8'h5c,8'h5c,8'h5e,8'h5f,8'h5e,8'h5e,8'h5c,8'h5b,8'h5f,8'h5d,8'h59,8'h58,8'h57,8'h44,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1a,8'h26,8'h2d,8'h39,8'h4a,8'h46,8'h24,8'h00,8'h00,8'h00,8'h0a,8'h48,8'h46,8'h3a,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'h12,8'h24,8'h2d,8'h31,8'h35,8'h39,8'h41,8'h40,8'h3d,8'h32,8'h22,8'h00,8'h00,8'h00,8'h00,8'h2a,8'h52,8'h5e,8'h5e,8'h58,8'h58,8'h29,8'h00,8'h00,8'h17,8'h47,8'h50,8'h4b,8'h49,8'h48,8'h48,8'h49,8'h44,8'h1e,8'h00,8'h00,8'h25,8'h55,8'h49,8'h43,8'h2f,8'h19,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h1b,8'h24,8'h30,8'h34,8'h40,8'h4c,8'h4e,8'h4d,8'h48,8'h44,8'h41,8'h40,8'h27,8'h5f,8'hdb,8'hd9,8'ha0,8'hbf,8'haa,8'hda,8'hb6,8'h4b,8'h63,8'h6f,8'h6a,8'h4c,8'h4a,8'h31,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h11,8'h25,8'h32,8'h35,8'h40,8'h48,8'h4e,8'h50,8'h43,8'h23,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h47,8'h58,8'h54,8'h57,8'h66,8'h74,8'h60,8'h6a,8'h5a,8'h4a,8'h41,8'h2b,8'h02,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h1f,8'h30,8'h3a,8'h47,8'h51,8'h4f,8'h51,8'h51,8'h52,8'h49,8'h38,8'h23,8'h0c,8'h00,8'h00,8'h0c,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h00,8'h00,8'h00,8'h25,8'h4c,8'h66,8'h64,8'h5f,8'h5e,8'h5d,8'h4f,8'h23,8'h00,8'h00,8'h00,8'h34,8'h5b,8'h59,8'h5a,8'h5e,8'h5e,8'h60,8'h62,8'h5f,8'h5b,8'h5a,8'h5a,8'h5b,8'h5b,8'h4b,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h13,8'h26,8'h42,8'h46,8'h4c,8'h4d,8'h4a,8'h2c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h12,8'h24,8'h2e,8'h3c,8'h47,8'h4b,8'h4c,8'h4b,8'h4d,8'h4e,8'h4b,8'h4e,8'h4d,8'h45,8'h25,8'h00,8'h00,8'h00,8'h00,8'h44,8'h5d,8'h5d,8'h5d,8'h5a,8'h25,8'h00,8'h00,8'h17,8'h44,8'h49,8'h48,8'h47,8'h46,8'h46,8'h48,8'h40,8'h15,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'h19,8'h26,8'h32,8'h41,8'h47,8'h4a,8'h4a,8'h4d,8'h4c,8'h4d,8'h50,8'h50,8'h4e,8'h4c,8'h42,8'h4e,8'hc9,8'hd2,8'h59,8'h2b,8'h79,8'h4b,8'h87,8'hbf,8'h5c,8'h81,8'h6d,8'h45,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h02,8'h16,8'h24,8'h33,8'h42,8'h45,8'h4c,8'h4c,8'h4c,8'h4f,8'h4f,8'h4d,8'h2c,8'h0c,8'h06,8'h11,8'h16,8'h0d,8'h00,8'h00,8'h00,8'h45,8'h53,8'h53,8'h57,8'h66,8'h7a,8'h51,8'h47,8'h29,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h1f,8'h28,8'h38,8'h49,8'h50,8'h56,8'h57,8'h54,8'h52,8'h52,8'h51,8'h54,8'h57,8'h58,8'h41,8'h1f,8'h00,8'h00,8'h00,8'h23,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h16,8'h00,8'h00,8'h10,8'h32,8'h5f,8'h64,8'h5d,8'h58,8'h57,8'h5c,8'h43,8'h03,8'h00,8'h00,8'h00,8'h4b,8'h5b,8'h58,8'h5c,8'h5e,8'h60,8'h62,8'h83,8'h6f,8'h5a,8'h5d,8'h5e,8'h55,8'h43,8'h21,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1c,8'h29,8'h3d,8'h47,8'h4f,8'h4a,8'h4a,8'h49,8'h3d,8'h16,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'h0e,8'h23,8'h2e,8'h3c,8'h45,8'h48,8'h4c,8'h4e,8'h4a,8'h49,8'h4c,8'h4d,8'h4f,8'h49,8'h47,8'h48,8'h4b,8'h42,8'h20,8'h00,8'h00,8'h00,8'h32,8'h53,8'h59,8'h64,8'h65,8'h27,8'h00,8'h00,8'h1e,8'h48,8'h4c,8'h4b,8'h4a,8'h49,8'h46,8'h49,8'h43,8'h1f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h05,8'h17,8'h24,8'h2f,8'h3f,8'h46,8'h4b,8'h4e,8'h4d,8'h4b,8'h4b,8'h4c,8'h4b,8'h4c,8'h4c,8'h4c,8'h49,8'h48,8'h42,8'h98,8'hbf,8'h53,8'h20,8'h00,8'h55,8'h42,8'h4b,8'hb6,8'h65,8'h62,8'h48,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h17,8'h23,8'h2b,8'h42,8'h4c,8'h4f,8'h4d,8'h4c,8'h4e,8'h4d,8'h49,8'h4b,8'h4e,8'h4d,8'h3a,8'h24,8'h2a,8'h36,8'h3d,8'h2b,8'h00,8'h00,8'h00,8'h46,8'h55,8'h52,8'h48,8'h39,8'h32,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h14,8'h25,8'h33,8'h45,8'h4b,8'h52,8'h54,8'h51,8'h53,8'h50,8'h4f,8'h4d,8'h50,8'h50,8'h55,8'h55,8'h58,8'h54,8'h2a,8'h10,8'h00,8'h00,8'h1f,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h23,8'h00,8'h00,8'h00,8'h28,8'h55,8'h61,8'h5f,8'h59,8'h56,8'h52,8'h4d,8'h28,8'h00,8'h00,8'h00,8'h2f,8'h5a,8'h5a,8'h5d,8'h5a,8'h68,8'h86,8'h67,8'h6d,8'h64,8'h5e,8'h61,8'h64,8'h57,8'h53,8'h51,8'h44,8'h00,8'h00,8'h00,8'h00,8'h0c,8'h23,8'h43,8'h49,8'h46,8'h4a,8'h4d,8'h49,8'h3f,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h02,8'h0c,8'h16,8'h27,8'h3b,8'h3a,8'h45,8'h4d,8'h4c,8'h49,8'h49,8'h49,8'h48,8'h47,8'h46,8'h47,8'h4b,8'h4b,8'h47,8'h47,8'h47,8'h48,8'h4b,8'h2f,8'h00,8'h00,8'h00,8'h2c,8'h5e,8'h5e,8'h6e,8'h69,8'h20,8'h00,8'h00,8'h24,8'h4c,8'h4d,8'h4a,8'h48,8'h48,8'h47,8'h49,8'h43,8'h17,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0f,8'h04,8'h0b,8'h20,8'h2f,8'h33,8'h3e,8'h48,8'h49,8'h49,8'h4b,8'h4c,8'h4b,8'h47,8'h45,8'h48,8'h48,8'h48,8'h49,8'h48,8'h46,8'h41,8'h6d,8'h86,8'h45,8'h15,8'h35,8'h00,8'h38,8'h45,8'h3e,8'h6f,8'h5c,8'h4a,8'h27,8'h00,8'h00,8'h00,8'h13,8'h28,8'h36,8'h42,8'h48,8'h4e,8'h4d,8'h4b,8'h4b,8'h4b,8'h4e,8'h48,8'h47,8'h4b,8'h4b,8'h4d,8'h4c,8'h46,8'h43,8'h44,8'h4d,8'h4f,8'h34,8'h00,8'h00,8'h00,8'h47,8'h43,8'h21,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h10,8'h26,8'h3d,8'h43,8'h49,8'h50,8'h53,8'h52,8'h51,8'h50,8'h4e,8'h51,8'h52,8'h4f,8'h52,8'h51,8'h51,8'h50,8'h52,8'h55,8'h57,8'h3a,8'h12,8'h00,8'h00,8'h0f,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h24,8'h00,8'h00,8'h00,8'h14,8'h42,8'h61,8'h5e,8'h59,8'h5a,8'h57,8'h56,8'h49,8'h1f,8'h00,8'h00,8'h00,8'h44,8'h5b,8'h59,8'h61,8'h6c,8'h6e,8'h86,8'h82,8'h67,8'h58,8'h63,8'h68,8'h5b,8'h5c,8'h6d,8'h77,8'h7b,8'h4d,8'h22,8'h00,8'h00,8'h00,8'h09,8'h3b,8'h4b,8'h46,8'h4b,8'h4a,8'h48,8'h2c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0b,8'h11,8'h0f,8'h13,8'h22,8'h25,8'h25,8'h26,8'h30,8'h47,8'h4a,8'h4a,8'h49,8'h46,8'h49,8'h46,8'h46,8'h47,8'h45,8'h45,8'h47,8'h49,8'h48,8'h4a,8'h3a,8'h00,8'h00,8'h00,8'h32,8'h83,8'h76,8'h82,8'h73,8'h13,8'h00,8'h00,8'h26,8'h4b,8'h48,8'h47,8'h45,8'h47,8'h49,8'h4b,8'h41,8'h08,8'h00,8'h00,8'h00,8'h00,8'h05,8'h0e,8'h0c,8'h09,8'h0c,8'h1a,8'h21,8'h21,8'h23,8'h2f,8'h43,8'h4b,8'h4d,8'h4a,8'h47,8'h45,8'h47,8'h48,8'h48,8'h4a,8'h4a,8'h3a,8'h45,8'h59,8'h38,8'h2a,8'h01,8'h2f,8'h00,8'h18,8'h3b,8'h46,8'h42,8'h45,8'h3d,8'h00,8'h00,8'h00,8'h18,8'h34,8'h48,8'h4d,8'h4a,8'h4b,8'h4c,8'h48,8'h45,8'h47,8'h45,8'h47,8'h46,8'h45,8'h4a,8'h47,8'h47,8'h49,8'h46,8'h45,8'h48,8'h4b,8'h4d,8'h31,8'h00,8'h00,8'h00,8'h46,8'h20,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0c,8'h09,8'h13,8'h23,8'h27,8'h29,8'h33,8'h42,8'h4c,8'h51,8'h52,8'h51,8'h52,8'h51,8'h4f,8'h50,8'h50,8'h4c,8'h4f,8'h50,8'h52,8'h56,8'h5a,8'h45,8'h14,8'h00,8'h00,8'h0b,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h1f,8'h00,8'h00,8'h01,8'h2a,8'h58,8'h63,8'h5b,8'h56,8'h58,8'h57,8'h55,8'h40,8'h03,8'h00,8'h00,8'h00,8'h4a,8'h5e,8'h5b,8'h68,8'h84,8'h69,8'h62,8'h75,8'h62,8'h6b,8'h77,8'h65,8'h5d,8'h69,8'h75,8'h75,8'h6e,8'h62,8'h4f,8'h2c,8'h00,8'h00,8'h00,8'h2c,8'h4b,8'h4a,8'h4b,8'h4c,8'h44,8'h1f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h11,8'h30,8'h4d,8'h4a,8'h49,8'h49,8'h48,8'h48,8'h48,8'h49,8'h49,8'h47,8'h49,8'h49,8'h48,8'h4a,8'h3c,8'h03,8'h00,8'h00,8'h35,8'h6d,8'h6b,8'h7f,8'h78,8'h18,8'h00,8'h00,8'h29,8'h4c,8'h48,8'h47,8'h48,8'h4b,8'h4a,8'h4d,8'h44,8'h10,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h11,8'h2f,8'h48,8'h46,8'h46,8'h47,8'h46,8'h49,8'h49,8'h49,8'h4a,8'h43,8'h24,8'h2b,8'h2e,8'h41,8'h35,8'h00,8'h00,8'h00,8'h06,8'h35,8'h59,8'h3d,8'h23,8'h17,8'h00,8'h00,8'h02,8'h2c,8'h49,8'h4a,8'h49,8'h4b,8'h4b,8'h49,8'h45,8'h46,8'h47,8'h45,8'h48,8'h43,8'h3c,8'h2f,8'h34,8'h47,8'h49,8'h47,8'h47,8'h49,8'h4a,8'h4a,8'h31,8'h00,8'h00,8'h01,8'h48,8'h30,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h10,8'h1e,8'h36,8'h4e,8'h52,8'h51,8'h4f,8'h4e,8'h4a,8'h4d,8'h4c,8'h50,8'h50,8'h4f,8'h54,8'h57,8'h5d,8'h4a,8'h20,8'h00,8'h00,8'h0b,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h25,8'h00,8'h00,8'h00,8'h21,8'h45,8'h64,8'h5d,8'h57,8'h55,8'h54,8'h55,8'h4d,8'h2d,8'h00,8'h00,8'h00,8'h27,8'h67,8'h6a,8'h5b,8'h6a,8'h6d,8'h68,8'h6f,8'h68,8'h5e,8'h6e,8'h6d,8'h5f,8'h67,8'h66,8'h6c,8'h70,8'h85,8'h65,8'h59,8'h4e,8'h16,8'h00,8'h00,8'h21,8'h41,8'h4d,8'h4c,8'h4c,8'h49,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h48,8'h4a,8'h48,8'h4d,8'h4a,8'h4a,8'h4b,8'h48,8'h49,8'h48,8'h46,8'h48,8'h47,8'h48,8'h39,8'h00,8'h00,8'h00,8'h39,8'h61,8'h57,8'h76,8'h71,8'h09,8'h00,8'h00,8'h2b,8'h49,8'h47,8'h48,8'h4a,8'h4b,8'h4b,8'h4d,8'h45,8'h12,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h24,8'h48,8'h49,8'h48,8'h48,8'h4a,8'h48,8'h47,8'h4b,8'h49,8'h27,8'h1e,8'h37,8'h45,8'h4a,8'h34,8'h00,8'h00,8'h00,8'h0f,8'h51,8'h7e,8'h4e,8'h1f,8'h00,8'h00,8'h00,8'h12,8'h40,8'h4b,8'h4c,8'h4b,8'h4e,8'h49,8'h45,8'h45,8'h46,8'h43,8'h3a,8'h2b,8'h1e,8'h17,8'h1b,8'h39,8'h4f,8'h4a,8'h48,8'h49,8'h4a,8'h4b,8'h48,8'h29,8'h00,8'h00,8'h10,8'h4d,8'h5a,8'h52,8'h51,8'h4e,8'h51,8'h42,8'h31,8'h27,8'h07,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h22,8'h47,8'h50,8'h4e,8'h4d,8'h4c,8'h4b,8'h4e,8'h51,8'h53,8'h51,8'h51,8'h52,8'h52,8'h5a,8'h4a,8'h22,8'h00,8'h00,8'h09,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h1e,8'h00,8'h00,8'h1a,8'h2a,8'h5a,8'h63,8'h5d,8'h5b,8'h57,8'h57,8'h57,8'h4b,8'h20,8'h00,8'h00,8'h00,8'h40,8'h7a,8'h81,8'h71,8'h6a,8'h6f,8'h6e,8'h6c,8'h65,8'h63,8'h6a,8'h62,8'h5c,8'h63,8'h67,8'h5d,8'h61,8'h6a,8'h5a,8'h57,8'h58,8'h34,8'h00,8'h00,8'h07,8'h35,8'h4a,8'h4c,8'h4b,8'h4a,8'h36,8'h00,8'h00,8'h00,8'h00,8'h22,8'h4b,8'h50,8'h4d,8'h34,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'h2b,8'h4b,8'h4c,8'h49,8'h4b,8'h49,8'h49,8'h49,8'h46,8'h46,8'h49,8'h46,8'h46,8'h45,8'h4b,8'h37,8'h00,8'h00,8'h00,8'h41,8'h65,8'h5f,8'h83,8'h6b,8'h00,8'h00,8'h00,8'h2c,8'h4a,8'h47,8'h47,8'h4a,8'h48,8'h49,8'h4a,8'h3f,8'h07,8'h00,8'h00,8'h1b,8'h26,8'h25,8'h24,8'h11,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0f,8'h2c,8'h47,8'h48,8'h48,8'h4b,8'h4d,8'h49,8'h49,8'h4a,8'h41,8'h27,8'h3f,8'h4a,8'h49,8'h47,8'h2a,8'h00,8'h00,8'h00,8'h23,8'h4d,8'h6e,8'h56,8'h30,8'h00,8'h00,8'h00,8'h20,8'h43,8'h4c,8'h48,8'h47,8'h48,8'h4b,8'h48,8'h42,8'h34,8'h24,8'h17,8'h01,8'h00,8'h01,8'h1f,8'h44,8'h4f,8'h4a,8'h48,8'h4a,8'h4a,8'h48,8'h43,8'h20,8'h00,8'h00,8'h23,8'h53,8'h7d,8'h74,8'h71,8'h63,8'h61,8'h57,8'h5d,8'h5e,8'h55,8'h54,8'h40,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h4b,8'h54,8'h52,8'h53,8'h52,8'h53,8'h56,8'h55,8'h53,8'h50,8'h51,8'h54,8'h52,8'h5b,8'h4c,8'h20,8'h00,8'h00,8'h0b,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h23,8'h00,8'h00,8'h00,8'h1b,8'h3c,8'h5e,8'h5d,8'h5a,8'h58,8'h57,8'h55,8'h53,8'h43,8'h08,8'h00,8'h00,8'h00,8'h4c,8'h61,8'h73,8'h83,8'h83,8'h7a,8'h65,8'h60,8'h6c,8'h69,8'h67,8'h60,8'h5b,8'h62,8'h65,8'h5d,8'h5f,8'h60,8'h55,8'h5f,8'h66,8'h38,8'h00,8'h00,8'h05,8'h36,8'h4e,8'h4b,8'h4d,8'h4c,8'h45,8'h1d,8'h00,8'h00,8'h00,8'h29,8'h6d,8'h78,8'h4f,8'h13,8'h00,8'h00,8'h00,8'h00,8'h00,8'h10,8'h26,8'h40,8'h4b,8'h4b,8'h49,8'h4d,8'h49,8'h47,8'h49,8'h48,8'h48,8'h49,8'h46,8'h45,8'h45,8'h48,8'h33,8'h00,8'h00,8'h00,8'h40,8'h71,8'h74,8'h6e,8'h59,8'h00,8'h00,8'h00,8'h2c,8'h4a,8'h47,8'h48,8'h4a,8'h47,8'h48,8'h49,8'h3e,8'h07,8'h00,8'h00,8'h21,8'h27,8'h26,8'h26,8'h26,8'h17,8'h00,8'h00,8'h00,8'h00,8'h11,8'h23,8'h43,8'h4b,8'h49,8'h49,8'h4a,8'h49,8'h4a,8'h48,8'h4a,8'h47,8'h46,8'h4e,8'h4e,8'h49,8'h48,8'h29,8'h00,8'h00,8'h00,8'h3a,8'h56,8'h5e,8'h56,8'h46,8'h00,8'h00,8'h00,8'h29,8'h48,8'h49,8'h49,8'h48,8'h46,8'h4b,8'h40,8'h27,8'h10,8'h00,8'h00,8'h00,8'h00,8'h02,8'h22,8'h46,8'h4d,8'h4c,8'h4b,8'h49,8'h49,8'h49,8'h3f,8'h11,8'h00,8'h00,8'h2b,8'h59,8'h6f,8'h6b,8'h61,8'h61,8'h5b,8'h56,8'h68,8'h7e,8'h6d,8'h66,8'h37,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0a,8'h33,8'h52,8'h54,8'h56,8'h58,8'h56,8'h57,8'h56,8'h51,8'h52,8'h50,8'h54,8'h58,8'h58,8'h5e,8'h48,8'h1f,8'h00,8'h00,8'h0d,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h1e,8'h00,8'h00,8'h00,8'h23,8'h4f,8'h60,8'h58,8'h56,8'h55,8'h53,8'h52,8'h52,8'h3f,8'h00,8'h00,8'h00,8'h00,8'h50,8'h5d,8'h5d,8'h6a,8'h87,8'h79,8'h5f,8'h63,8'h89,8'h6d,8'h5b,8'h59,8'h5a,8'h5b,8'h5f,8'h60,8'h60,8'h6c,8'h6e,8'h87,8'h68,8'h27,8'h00,8'h00,8'h0c,8'h3a,8'h54,8'h50,8'h4d,8'h4c,8'h4a,8'h2c,8'h00,8'h00,8'h00,8'h00,8'h69,8'h6b,8'h3d,8'h00,8'h00,8'h00,8'h00,8'h0c,8'h25,8'h37,8'h45,8'h48,8'h48,8'h46,8'h45,8'h48,8'h48,8'h47,8'h42,8'h41,8'h48,8'h47,8'h47,8'h48,8'h48,8'h48,8'h32,8'h00,8'h00,8'h00,8'h4e,8'h8d,8'h7b,8'h7a,8'h59,8'h00,8'h00,8'h00,8'h2c,8'h48,8'h46,8'h47,8'h49,8'h47,8'h46,8'h49,8'h42,8'h09,8'h00,8'h00,8'h22,8'h26,8'h26,8'h26,8'h24,8'h00,8'h00,8'h00,8'h14,8'h1f,8'h2b,8'h44,8'h48,8'h4b,8'h4b,8'h47,8'h47,8'h44,8'h36,8'h2d,8'h46,8'h4b,8'h49,8'h49,8'h47,8'h48,8'h47,8'h28,8'h00,8'h00,8'h00,8'h44,8'h62,8'h5e,8'h5b,8'h45,8'h00,8'h00,8'h05,8'h31,8'h48,8'h48,8'h4b,8'h49,8'h45,8'h36,8'h1d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h09,8'h28,8'h4a,8'h4e,8'h50,8'h4a,8'h49,8'h4b,8'h4c,8'h33,8'h03,8'h00,8'h00,8'h39,8'h5c,8'h5a,8'h5a,8'h5d,8'h60,8'h60,8'h61,8'h6a,8'h87,8'h6e,8'h49,8'h00,8'h00,8'h00,8'h00,8'h10,8'h13,8'h2c,8'h49,8'h4d,8'h4c,8'h50,8'h52,8'h50,8'h4d,8'h3a,8'h2d,8'h4b,8'h4e,8'h4e,8'h50,8'h50,8'h57,8'h44,8'h14,8'h00,8'h00,8'h0b,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h26,8'h06,8'h00,8'h00,8'h13,8'h31,8'h5e,8'h5a,8'h59,8'h55,8'h56,8'h55,8'h51,8'h54,8'h37,8'h00,8'h00,8'h00,8'h1b,8'h5b,8'h75,8'h71,8'h64,8'h78,8'h63,8'h5b,8'h5d,8'h6b,8'h5f,8'h5c,8'h59,8'h58,8'h58,8'h5e,8'h64,8'h6a,8'h85,8'h7b,8'h85,8'h55,8'h00,8'h00,8'h00,8'h22,8'h43,8'h4f,8'h4c,8'h4c,8'h4c,8'h4c,8'h3f,8'h09,8'h00,8'h00,8'h00,8'h3f,8'h69,8'h44,8'h00,8'h00,8'h00,8'h18,8'h3a,8'h47,8'h4a,8'h48,8'h46,8'h48,8'h47,8'h46,8'h45,8'h44,8'h33,8'h1f,8'h29,8'h49,8'h45,8'h44,8'h45,8'h45,8'h47,8'h34,8'h00,8'h00,8'h00,8'h4a,8'h94,8'h83,8'h8c,8'h5b,8'h00,8'h00,8'h00,8'h29,8'h48,8'h45,8'h45,8'h46,8'h44,8'h41,8'h43,8'h3d,8'h03,8'h00,8'h00,8'h21,8'h26,8'h26,8'h26,8'h15,8'h00,8'h00,8'h16,8'h22,8'h36,8'h41,8'h42,8'h44,8'h46,8'h44,8'h42,8'h3a,8'h24,8'h16,8'h1f,8'h33,8'h3f,8'h3c,8'h3b,8'h39,8'h39,8'h38,8'h22,8'h00,8'h00,8'h00,8'h55,8'h6f,8'h5c,8'h6a,8'h44,8'h00,8'h00,8'h0b,8'h28,8'h34,8'h33,8'h33,8'h33,8'h31,8'h1d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h07,8'h25,8'h34,8'h2f,8'h2f,8'h2f,8'h30,8'h31,8'h32,8'h24,8'h00,8'h00,8'h00,8'h43,8'h5c,8'h5e,8'h59,8'h5c,8'h64,8'h6a,8'h6e,8'h67,8'h7c,8'h62,8'h28,8'h00,8'h00,8'h02,8'h13,8'h16,8'h1a,8'h27,8'h27,8'h27,8'h26,8'h28,8'h28,8'h29,8'h25,8'h20,8'h1f,8'h27,8'h28,8'h26,8'h26,8'h27,8'h29,8'h24,8'h0f,8'h00,8'h00,8'h09,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h26,8'h23,8'h00,8'h00,8'h00,8'h1d,8'h3d,8'h4d,8'h4c,8'h4a,8'h45,8'h45,8'h44,8'h46,8'h47,8'h25,8'h00,8'h00,8'h00,8'h2e,8'h69,8'h78,8'h7c,8'h5c,8'h60,8'h58,8'h59,8'h5c,8'h5e,8'h60,8'h5e,8'h5a,8'h59,8'h59,8'h60,8'h6f,8'h74,8'h68,8'h58,8'h47,8'h14,8'h00,8'h00,8'h09,8'h22,8'h31,8'h3a,8'h3a,8'h36,8'h34,8'h34,8'h2c,8'h13,8'h00,8'h00,8'h00,8'h29,8'h6b,8'h3e,8'h00,8'h00,8'h0b,8'h20,8'h31,8'h2e,8'h2e,8'h2c,8'h2a,8'h2b,8'h2d,8'h2b,8'h28,8'h23,8'h11,8'h0a,8'h1b,8'h2b,8'h2b,8'h2a,8'h2a,8'h29,8'h29,8'h23,8'h00,8'h00,8'h00,8'h4d,8'h72,8'h6e,8'h66,8'h4f,8'h00,8'h00,8'h00,8'h18,8'h26,8'h27,8'h28,8'h27,8'h26,8'h27,8'h25,8'h20,8'h00,8'h00,8'h00,8'h21,8'h26,8'h26,8'h26,8'h00,8'h00,8'h10,8'h18,8'h1f,8'h23,8'h23,8'h23,8'h23,8'h21,8'h18,8'h15,8'h14,8'h00,8'h00,8'h13,8'h20,8'h23,8'h20,8'h20,8'h20,8'h1f,8'h1a,8'h0f,8'h00,8'h00,8'h09,8'h74,8'h7d,8'h5d,8'h5f,8'h34,8'h00,8'h00,8'h0c,8'h15,8'h1a,8'h1d,8'h1d,8'h19,8'h18,8'h0c,8'h00,8'h00,8'h00,8'h0e,8'h00,8'h00,8'h00,8'h12,8'h20,8'h1f,8'h21,8'h21,8'h22,8'h1f,8'h19,8'h13,8'h0d,8'h00,8'h00,8'h23,8'h50,8'h59,8'h5c,8'h5b,8'h64,8'h6b,8'h6a,8'h6d,8'h63,8'h6a,8'h52,8'h00,8'h00,8'h00,8'h18,8'h1f,8'h20,8'h21,8'h21,8'h21,8'h21,8'h22,8'h1e,8'h0d,8'h0a,8'h00,8'h1a,8'h13,8'h20,8'h23,8'h23,8'h23,8'h24,8'h23,8'h1f,8'h0c,8'h00,8'h00,8'h0d,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h18,8'h00,8'h00,8'h15,8'h12,8'h20,8'h23,8'h26,8'h25,8'h23,8'h22,8'h24,8'h26,8'h22,8'h15,8'h00,8'h00,8'h00,8'h44,8'h75,8'h5e,8'h5a,8'h58,8'h5d,8'h5b,8'h5b,8'h58,8'h59,8'h5d,8'h5a,8'h59,8'h60,8'h67,8'h7b,8'h81,8'h81,8'h62,8'h34,8'h00,8'h00,8'h00,8'h04,8'h1f,8'h24,8'h27,8'h27,8'h27,8'h27,8'h26,8'h24,8'h24,8'h20,8'h02,8'h00,8'h00,8'h00,8'h44,8'h2b,8'h00,8'h00,8'h13,8'h1d,8'h23,8'h23,8'h26,8'h27,8'h25,8'h21,8'h15,8'h03,8'h00,8'h00,8'h00,8'h0e,8'h16,8'h26,8'h27,8'h27,8'h27,8'h24,8'h23,8'h20,8'h00,8'h00,8'h00,8'h64,8'h6e,8'h57,8'h65,8'h53,8'h00,8'h00,8'h00,8'h19,8'h27,8'h29,8'h2c,8'h2b,8'h2a,8'h2a,8'h2a,8'h22,8'h00,8'h00,8'h00,8'h21,8'h26,8'h26,8'h25,8'h00,8'h00,8'h13,8'h23,8'h27,8'h28,8'h2a,8'h29,8'h29,8'h21,8'h0b,8'h00,8'h00,8'h00,8'h00,8'h17,8'h29,8'h2d,8'h2e,8'h2d,8'h2d,8'h2d,8'h29,8'h16,8'h00,8'h00,8'h11,8'h6c,8'h7c,8'h69,8'h55,8'h1a,8'h00,8'h00,8'h10,8'h27,8'h2e,8'h2e,8'h30,8'h2d,8'h1f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h15,8'h20,8'h2a,8'h2f,8'h31,8'h30,8'h32,8'h2e,8'h2a,8'h1c,8'h00,8'h00,8'h00,8'h37,8'h59,8'h5c,8'h5f,8'h5f,8'h62,8'h63,8'h67,8'h67,8'h5f,8'h75,8'h54,8'h00,8'h00,8'h01,8'h1b,8'h27,8'h2c,8'h31,8'h32,8'h31,8'h2a,8'h22,8'h18,8'h00,8'h00,8'h00,8'h08,8'h1f,8'h2f,8'h34,8'h36,8'h34,8'h36,8'h30,8'h23,8'h0d,8'h00,8'h00,8'h0a,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h00,8'h00},
'{8'h00,8'h00,8'h26,8'h25,8'h00,8'h00,8'h00,8'h17,8'h1f,8'h26,8'h2a,8'h2a,8'h2b,8'h2d,8'h2f,8'h2f,8'h2d,8'h28,8'h16,8'h00,8'h00,8'h00,8'h33,8'h62,8'h59,8'h5a,8'h5c,8'h5c,8'h5e,8'h5c,8'h5a,8'h58,8'h64,8'h6c,8'h61,8'h6a,8'h71,8'h87,8'h69,8'h5c,8'h2b,8'h00,8'h00,8'h00,8'h03,8'h12,8'h23,8'h2e,8'h34,8'h31,8'h33,8'h32,8'h31,8'h2d,8'h2e,8'h27,8'h10,8'h00,8'h00,8'h00,8'h1b,8'h00,8'h00,8'h00,8'h14,8'h24,8'h2d,8'h2e,8'h2f,8'h2c,8'h2d,8'h24,8'h0d,8'h00,8'h00,8'h00,8'h00,8'h0c,8'h22,8'h2c,8'h2f,8'h30,8'h31,8'h2c,8'h29,8'h1f,8'h00,8'h00,8'h00,8'h61,8'h73,8'h60,8'h67,8'h49,8'h00,8'h00,8'h00,8'h1f,8'h2b,8'h2e,8'h30,8'h2f,8'h2f,8'h2e,8'h2e,8'h25,8'h00,8'h00,8'h00,8'h21,8'h27,8'h26,8'h24,8'h00,8'h00,8'h18,8'h28,8'h2a,8'h2d,8'h30,8'h2d,8'h2a,8'h14,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1b,8'h2a,8'h31,8'h32,8'h31,8'h31,8'h31,8'h2b,8'h14,8'h00,8'h00,8'h24,8'h5c,8'h7b,8'h6b,8'h46,8'h00,8'h00,8'h02,8'h19,8'h2c,8'h30,8'h30,8'h2f,8'h30,8'h1f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'h15,8'h18,8'h26,8'h2e,8'h2f,8'h32,8'h2c,8'h2c,8'h2b,8'h29,8'h13,8'h00,8'h00,8'h00,8'h55,8'h59,8'h5e,8'h60,8'h64,8'h69,8'h5d,8'h63,8'h7f,8'h63,8'h60,8'h3c,8'h00,8'h00,8'h07,8'h1f,8'h2a,8'h2f,8'h35,8'h35,8'h2f,8'h24,8'h0d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1f,8'h30,8'h34,8'h36,8'h35,8'h36,8'h31,8'h23,8'h10,8'h00,8'h00,8'h0c,8'h26,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h24,8'h23,8'h16,8'h20,8'h26,8'h00},
'{8'h00,8'h00,8'h26,8'h20,8'h00,8'h00,8'h18,8'h1e,8'h23,8'h27,8'h2c,8'h2e,8'h31,8'h35,8'h37,8'h33,8'h30,8'h2b,8'h1a,8'h00,8'h00,8'h00,8'h15,8'h4f,8'h5a,8'h5a,8'h58,8'h58,8'h5c,8'h5d,8'h5b,8'h5a,8'h69,8'h7c,8'h6a,8'h6f,8'h65,8'h58,8'h3c,8'h15,8'h00,8'h00,8'h00,8'h13,8'h23,8'h24,8'h2e,8'h35,8'h36,8'h35,8'h33,8'h33,8'h30,8'h30,8'h30,8'h2d,8'h22,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1c,8'h27,8'h2e,8'h2e,8'h30,8'h2b,8'h2a,8'h21,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0b,8'h23,8'h29,8'h2d,8'h31,8'h30,8'h2d,8'h29,8'h14,8'h00,8'h00,8'h00,8'h63,8'h5e,8'h49,8'h41,8'h20,8'h00,8'h00,8'h00,8'h1f,8'h2a,8'h2c,8'h2f,8'h2f,8'h2f,8'h31,8'h2e,8'h25,8'h00,8'h00,8'h00,8'h21,8'h27,8'h26,8'h1f,8'h00,8'h00,8'h1f,8'h2b,8'h2c,8'h2e,8'h30,8'h2e,8'h26,8'h0b,8'h00,8'h00,8'h04,8'h00,8'h00,8'h1d,8'h2a,8'h32,8'h32,8'h31,8'h30,8'h2f,8'h27,8'h0a,8'h00,8'h00,8'h23,8'h51,8'h62,8'h4f,8'h1d,8'h00,8'h00,8'h08,8'h1e,8'h2a,8'h2f,8'h32,8'h31,8'h2f,8'h1c,8'h07,8'h07,8'h0a,8'h1c,8'h21,8'h21,8'h24,8'h28,8'h2b,8'h2b,8'h2e,8'h2e,8'h27,8'h24,8'h20,8'h11,8'h00,8'h00,8'h00,8'h3f,8'h6f,8'h67,8'h66,8'h63,8'h63,8'h66,8'h60,8'h65,8'h74,8'h67,8'h5b,8'h28,8'h00,8'h00,8'h0e,8'h21,8'h2d,8'h33,8'h34,8'h31,8'h2f,8'h22,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1f,8'h33,8'h35,8'h34,8'h35,8'h33,8'h30,8'h24,8'h19,8'h00,8'h00,8'h0b,8'h26,8'h00,8'h24,8'h22,8'h20,8'h1e,8'h09,8'h00,8'h00,8'h00,8'h11,8'h26,8'h26},
'{8'h00,8'h26,8'h26,8'h09,8'h00,8'h00,8'h13,8'h1e,8'h26,8'h27,8'h2c,8'h2f,8'h34,8'h35,8'h33,8'h31,8'h33,8'h30,8'h23,8'h00,8'h00,8'h00,8'h00,8'h39,8'h50,8'h59,8'h57,8'h56,8'h58,8'h5b,8'h5b,8'h5c,8'h62,8'h5a,8'h66,8'h64,8'h3e,8'h0f,8'h00,8'h00,8'h00,8'h00,8'h20,8'h29,8'h2f,8'h33,8'h37,8'h37,8'h36,8'h34,8'h33,8'h33,8'h32,8'h32,8'h31,8'h2d,8'h28,8'h19,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1f,8'h29,8'h2e,8'h2e,8'h30,8'h2b,8'h28,8'h1c,8'h00,8'h00,8'h10,8'h00,8'h00,8'h16,8'h27,8'h2a,8'h2f,8'h30,8'h2f,8'h2d,8'h2c,8'h18,8'h00,8'h00,8'h00,8'h32,8'h2e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h2b,8'h2c,8'h31,8'h32,8'h33,8'h33,8'h2f,8'h25,8'h00,8'h00,8'h00,8'h21,8'h27,8'h27,8'h11,8'h00,8'h0a,8'h20,8'h2b,8'h2f,8'h33,8'h31,8'h2f,8'h26,8'h00,8'h00,8'h00,8'h22,8'h00,8'h00,8'h1f,8'h2c,8'h34,8'h34,8'h33,8'h30,8'h2d,8'h22,8'h05,8'h00,8'h00,8'h23,8'h44,8'h2d,8'h00,8'h00,8'h00,8'h00,8'h0c,8'h21,8'h2c,8'h2e,8'h32,8'h32,8'h31,8'h24,8'h1f,8'h23,8'h25,8'h2a,8'h2c,8'h2c,8'h31,8'h30,8'h2c,8'h2b,8'h2a,8'h25,8'h16,8'h0c,8'h00,8'h00,8'h00,8'h00,8'h26,8'h5a,8'h63,8'h85,8'h76,8'h5f,8'h5f,8'h5d,8'h67,8'h7a,8'h6e,8'h79,8'h63,8'h17,8'h00,8'h00,8'h17,8'h24,8'h31,8'h36,8'h32,8'h2f,8'h2d,8'h23,8'h00,8'h00,8'h10,8'h0c,8'h00,8'h04,8'h20,8'h33,8'h38,8'h37,8'h35,8'h33,8'h33,8'h23,8'h1d,8'h00,8'h00,8'h00,8'h21,8'h0e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h26,8'h00},
'{8'h00,8'h26,8'h24,8'h00,8'h00,8'h00,8'h14,8'h1f,8'h2a,8'h2b,8'h30,8'h34,8'h38,8'h38,8'h35,8'h34,8'h37,8'h35,8'h25,8'h0b,8'h00,8'h00,8'h00,8'h00,8'h2d,8'h47,8'h4a,8'h4c,8'h50,8'h54,8'h54,8'h51,8'h4e,8'h47,8'h41,8'h21,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h34,8'h32,8'h33,8'h37,8'h36,8'h35,8'h35,8'h35,8'h35,8'h35,8'h34,8'h32,8'h30,8'h2e,8'h2c,8'h23,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1e,8'h2a,8'h30,8'h31,8'h2f,8'h2c,8'h28,8'h11,8'h00,8'h00,8'h1f,8'h00,8'h00,8'h1f,8'h2a,8'h2e,8'h30,8'h31,8'h30,8'h2e,8'h2d,8'h1c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h08,8'h21,8'h2b,8'h2e,8'h33,8'h33,8'h32,8'h2f,8'h2f,8'h27,8'h00,8'h00,8'h00,8'h21,8'h27,8'h27,8'h09,8'h00,8'h12,8'h24,8'h30,8'h34,8'h31,8'h2f,8'h2c,8'h21,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h22,8'h2f,8'h32,8'h32,8'h34,8'h31,8'h2f,8'h23,8'h02,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0c,8'h24,8'h2f,8'h31,8'h34,8'h34,8'h34,8'h2f,8'h2e,8'h30,8'h2e,8'h2d,8'h2f,8'h2f,8'h30,8'h2f,8'h2c,8'h26,8'h23,8'h15,8'h00,8'h00,8'h00,8'h00,8'h00,8'h36,8'h56,8'h5d,8'h60,8'h69,8'h63,8'h5c,8'h5a,8'h59,8'h65,8'h74,8'h80,8'ha3,8'h68,8'h00,8'h00,8'h00,8'h14,8'h27,8'h33,8'h33,8'h35,8'h30,8'h29,8'h1f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h10,8'h21,8'h34,8'h38,8'h3a,8'h37,8'h35,8'h32,8'h24,8'h12,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h00,8'h00,8'h00},
'{8'h00,8'h26,8'h15,8'h00,8'h00,8'h11,8'h1a,8'h26,8'h2c,8'h2c,8'h30,8'h35,8'h36,8'h38,8'h38,8'h37,8'h33,8'h33,8'h2d,8'h1f,8'h03,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1b,8'h20,8'h22,8'h22,8'h1e,8'h13,8'h00,8'h00,8'h00,8'h00,8'h00,8'h05,8'h1f,8'h27,8'h2e,8'h35,8'h3a,8'h3a,8'h36,8'h35,8'h36,8'h36,8'h34,8'h36,8'h35,8'h33,8'h31,8'h30,8'h32,8'h30,8'h27,8'h0a,8'h00,8'h00,8'h00,8'h00,8'h09,8'h1f,8'h2c,8'h2e,8'h30,8'h2f,8'h2c,8'h26,8'h05,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1f,8'h2d,8'h33,8'h33,8'h33,8'h31,8'h2d,8'h2b,8'h19,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0a,8'h21,8'h2a,8'h2e,8'h33,8'h31,8'h32,8'h32,8'h30,8'h27,8'h00,8'h00,8'h00,8'h22,8'h27,8'h25,8'h00,8'h00,8'h18,8'h29,8'h32,8'h35,8'h32,8'h30,8'h2c,8'h1f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h17,8'h28,8'h33,8'h33,8'h32,8'h34,8'h32,8'h31,8'h23,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h13,8'h25,8'h2f,8'h32,8'h33,8'h34,8'h34,8'h32,8'h30,8'h30,8'h32,8'h30,8'h2f,8'h30,8'h30,8'h2b,8'h21,8'h07,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2c,8'h51,8'h62,8'h67,8'h5d,8'h5b,8'h5a,8'h5a,8'h5b,8'h5b,8'h61,8'h6f,8'h75,8'h87,8'h87,8'h58,8'h00,8'h00,8'h00,8'h1f,8'h2c,8'h33,8'h34,8'h34,8'h30,8'h28,8'h16,8'h00,8'h00,8'h00,8'h00,8'h00,8'h13,8'h26,8'h32,8'h38,8'h36,8'h36,8'h36,8'h32,8'h20,8'h0a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h01,8'h14,8'h1f,8'h00,8'h00,8'h00,8'h25,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h25,8'h00,8'h00,8'h00,8'h19,8'h19,8'h29,8'h2d,8'h2f,8'h31,8'h33,8'h35,8'h38,8'h38,8'h38,8'h36,8'h34,8'h32,8'h28,8'h1b,8'h0a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h1a,8'h1f,8'h27,8'h31,8'h33,8'h3a,8'h37,8'h3a,8'h37,8'h38,8'h39,8'h37,8'h34,8'h35,8'h35,8'h35,8'h31,8'h31,8'h34,8'h31,8'h2d,8'h20,8'h00,8'h00,8'h00,8'h00,8'h10,8'h20,8'h2d,8'h2f,8'h30,8'h30,8'h2b,8'h23,8'h00,8'h00,8'h00,8'h00,8'h00,8'h10,8'h20,8'h2e,8'h32,8'h32,8'h35,8'h33,8'h2e,8'h2b,8'h18,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h09,8'h05,8'h00,8'h00,8'h12,8'h24,8'h2b,8'h2c,8'h32,8'h31,8'h32,8'h31,8'h30,8'h26,8'h00,8'h00,8'h00,8'h22,8'h27,8'h25,8'h00,8'h00,8'h20,8'h2a,8'h32,8'h33,8'h34,8'h30,8'h2c,8'h1e,8'h00,8'h00,8'h00,8'h00,8'h15,8'h23,8'h2a,8'h30,8'h34,8'h33,8'h35,8'h32,8'h31,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'h0d,8'h00,8'h00,8'h17,8'h26,8'h2d,8'h31,8'h2f,8'h2f,8'h30,8'h30,8'h31,8'h32,8'h32,8'h2e,8'h2d,8'h2f,8'h2c,8'h23,8'h05,8'h00,8'h00,8'h00,8'h00,8'h27,8'h46,8'h6b,8'h84,8'h66,8'h69,8'h67,8'h5a,8'h56,8'h58,8'h5d,8'h5b,8'h62,8'h82,8'h8b,8'h8e,8'h84,8'h44,8'h00,8'h00,8'h03,8'h21,8'h2d,8'h32,8'h35,8'h33,8'h35,8'h29,8'h0a,8'h00,8'h00,8'h00,8'h05,8'h14,8'h21,8'h29,8'h2d,8'h35,8'h34,8'h35,8'h33,8'h2e,8'h1f,8'h0f,8'h00,8'h00,8'h00,8'h0c,8'h12,8'h14,8'h17,8'h00,8'h00,8'h00,8'h25,8'h26,8'h00,8'h00,8'h00,8'h00},
'{8'h26,8'h25,8'h00,8'h00,8'h00,8'h10,8'h1b,8'h29,8'h2d,8'h2f,8'h33,8'h34,8'h36,8'h37,8'h3a,8'h3a,8'h3a,8'h38,8'h37,8'h34,8'h2a,8'h1d,8'h18,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h09,8'h1c,8'h1c,8'h24,8'h2a,8'h31,8'h33,8'h37,8'h39,8'h38,8'h3a,8'h39,8'h39,8'h3b,8'h39,8'h38,8'h35,8'h35,8'h34,8'h34,8'h32,8'h31,8'h2e,8'h2c,8'h25,8'h0b,8'h00,8'h00,8'h00,8'h10,8'h23,8'h2f,8'h2f,8'h2f,8'h33,8'h30,8'h23,8'h00,8'h00,8'h00,8'h00,8'h0a,8'h20,8'h29,8'h2f,8'h2f,8'h32,8'h35,8'h32,8'h2e,8'h2d,8'h18,8'h00,8'h00,8'h00,8'h05,8'h09,8'h0d,8'h0a,8'h00,8'h00,8'h00,8'h0d,8'h23,8'h2d,8'h2e,8'h32,8'h33,8'h31,8'h31,8'h2f,8'h26,8'h05,8'h00,8'h00,8'h22,8'h28,8'h21,8'h00,8'h00,8'h20,8'h2b,8'h31,8'h33,8'h33,8'h2e,8'h2b,8'h1f,8'h00,8'h00,8'h0e,8'h19,8'h22,8'h28,8'h2f,8'h32,8'h36,8'h34,8'h33,8'h34,8'h32,8'h25,8'h0b,8'h00,8'h00,8'h00,8'h06,8'h0d,8'h10,8'h0b,8'h00,8'h05,8'h14,8'h27,8'h2b,8'h2d,8'h2c,8'h2c,8'h2d,8'h2e,8'h2a,8'h27,8'h25,8'h22,8'h25,8'h2a,8'h27,8'h17,8'h00,8'h00,8'h00,8'h1e,8'h37,8'h50,8'h61,8'h6d,8'h7d,8'h67,8'h76,8'h58,8'h55,8'h59,8'h63,8'h5f,8'h58,8'h5a,8'h65,8'h83,8'h7d,8'h77,8'h36,8'h00,8'h00,8'h10,8'h21,8'h2d,8'h31,8'h33,8'h33,8'h30,8'h25,8'h11,8'h00,8'h00,8'h18,8'h19,8'h24,8'h2c,8'h32,8'h32,8'h32,8'h34,8'h37,8'h35,8'h2e,8'h21,8'h1d,8'h07,8'h0f,8'h1f,8'h12,8'h13,8'h21,8'h02,8'h00,8'h00,8'h21,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h26,8'h24,8'h00,8'h00,8'h00,8'h15,8'h1c,8'h29,8'h2d,8'h30,8'h32,8'h35,8'h37,8'h39,8'h3b,8'h3d,8'h3c,8'h3a,8'h38,8'h35,8'h34,8'h2d,8'h28,8'h26,8'h20,8'h0e,8'h06,8'h02,8'h08,8'h10,8'h14,8'h19,8'h1f,8'h23,8'h26,8'h2d,8'h2c,8'h2d,8'h32,8'h34,8'h34,8'h36,8'h36,8'h38,8'h39,8'h38,8'h39,8'h3a,8'h3b,8'h39,8'h37,8'h37,8'h35,8'h35,8'h33,8'h31,8'h2e,8'h2e,8'h2b,8'h18,8'h00,8'h00,8'h00,8'h14,8'h27,8'h2e,8'h30,8'h30,8'h30,8'h31,8'h2b,8'h1b,8'h11,8'h17,8'h20,8'h24,8'h2c,8'h30,8'h31,8'h2f,8'h31,8'h32,8'h32,8'h30,8'h2e,8'h24,8'h16,8'h11,8'h12,8'h15,8'h13,8'h03,8'h00,8'h00,8'h00,8'h00,8'h09,8'h21,8'h2d,8'h2e,8'h32,8'h33,8'h31,8'h31,8'h2e,8'h25,8'h01,8'h00,8'h00,8'h21,8'h28,8'h1f,8'h00,8'h0d,8'h24,8'h2e,8'h31,8'h33,8'h30,8'h2f,8'h31,8'h25,8'h12,8'h20,8'h26,8'h2c,8'h2c,8'h2f,8'h32,8'h34,8'h39,8'h36,8'h32,8'h31,8'h33,8'h2b,8'h14,8'h0f,8'h11,8'h1f,8'h1a,8'h0e,8'h00,8'h00,8'h00,8'h0c,8'h1e,8'h2a,8'h2c,8'h2e,8'h2d,8'h2d,8'h29,8'h22,8'h1e,8'h1a,8'h07,8'h0c,8'h15,8'h26,8'h21,8'h04,8'h00,8'h00,8'h00,8'h2d,8'h30,8'h2d,8'h29,8'h23,8'h25,8'h2a,8'h31,8'h2c,8'h33,8'h45,8'h81,8'h6e,8'h5b,8'h71,8'h6d,8'h68,8'h5e,8'h53,8'h24,8'h00,8'h00,8'h16,8'h26,8'h2e,8'h32,8'h35,8'h34,8'h30,8'h28,8'h15,8'h19,8'h21,8'h27,8'h2c,8'h2e,8'h30,8'h36,8'h36,8'h34,8'h36,8'h37,8'h35,8'h30,8'h24,8'h17,8'h12,8'h1d,8'h1e,8'h14,8'h0f,8'h00,8'h00,8'h00,8'h22,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h26,8'h24,8'h00,8'h00,8'h00,8'h18,8'h1f,8'h29,8'h2c,8'h33,8'h34,8'h35,8'h36,8'h38,8'h39,8'h3a,8'h3c,8'h3b,8'h38,8'h36,8'h34,8'h31,8'h2f,8'h2f,8'h2b,8'h26,8'h24,8'h25,8'h25,8'h24,8'h25,8'h26,8'h28,8'h2b,8'h2c,8'h2f,8'h31,8'h34,8'h36,8'h32,8'h33,8'h35,8'h37,8'h37,8'h39,8'h3a,8'h3a,8'h3a,8'h3b,8'h39,8'h3c,8'h39,8'h35,8'h34,8'h33,8'h2f,8'h2e,8'h32,8'h2a,8'h1e,8'h06,8'h00,8'h01,8'h1d,8'h29,8'h30,8'h32,8'h32,8'h31,8'h34,8'h35,8'h2e,8'h26,8'h27,8'h2c,8'h2c,8'h2f,8'h32,8'h31,8'h2e,8'h31,8'h30,8'h2f,8'h2e,8'h2e,8'h2b,8'h25,8'h21,8'h23,8'h1d,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0c,8'h24,8'h2c,8'h2b,8'h2f,8'h31,8'h2f,8'h30,8'h2d,8'h24,8'h00,8'h00,8'h00,8'h21,8'h27,8'h12,8'h00,8'h13,8'h27,8'h30,8'h31,8'h31,8'h30,8'h31,8'h37,8'h30,8'h27,8'h2b,8'h2f,8'h30,8'h2d,8'h2d,8'h33,8'h34,8'h35,8'h34,8'h30,8'h30,8'h31,8'h2d,8'h24,8'h1d,8'h21,8'h24,8'h1f,8'h00,8'h00,8'h00,8'h00,8'h14,8'h21,8'h29,8'h29,8'h26,8'h22,8'h1e,8'h11,8'h10,8'h00,8'h00,8'h00,8'h16,8'h21,8'h28,8'h19,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h2b,8'h31,8'h58,8'h83,8'h74,8'h67,8'h5e,8'h4f,8'h07,8'h00,8'h00,8'h14,8'h2a,8'h32,8'h32,8'h37,8'h36,8'h32,8'h2f,8'h27,8'h25,8'h2d,8'h33,8'h32,8'h32,8'h33,8'h34,8'h33,8'h35,8'h32,8'h30,8'h32,8'h31,8'h2c,8'h26,8'h27,8'h24,8'h1c,8'h18,8'h00,8'h00,8'h00,8'h22,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h26,8'h24,8'h00,8'h00,8'h00,8'h13,8'h20,8'h2a,8'h2c,8'h31,8'h33,8'h35,8'h37,8'h36,8'h38,8'h39,8'h39,8'h3a,8'h38,8'h39,8'h36,8'h34,8'h34,8'h35,8'h33,8'h30,8'h2f,8'h2f,8'h2f,8'h2d,8'h2e,8'h30,8'h30,8'h30,8'h2e,8'h30,8'h32,8'h35,8'h36,8'h35,8'h36,8'h37,8'h39,8'h39,8'h37,8'h39,8'h3a,8'h3b,8'h3a,8'h38,8'h37,8'h35,8'h37,8'h38,8'h33,8'h2d,8'h29,8'h25,8'h20,8'h14,8'h00,8'h00,8'h0a,8'h1a,8'h2b,8'h30,8'h33,8'h34,8'h38,8'h37,8'h34,8'h35,8'h33,8'h33,8'h31,8'h2f,8'h30,8'h33,8'h32,8'h2e,8'h2f,8'h2f,8'h2f,8'h2f,8'h2e,8'h2d,8'h2d,8'h26,8'h1d,8'h02,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0a,8'h24,8'h2e,8'h2f,8'h32,8'h30,8'h35,8'h31,8'h2e,8'h25,8'h01,8'h00,8'h00,8'h22,8'h25,8'h00,8'h00,8'h14,8'h2a,8'h31,8'h31,8'h32,8'h32,8'h34,8'h35,8'h32,8'h31,8'h30,8'h31,8'h31,8'h2e,8'h2e,8'h31,8'h31,8'h32,8'h31,8'h30,8'h2f,8'h30,8'h2f,8'h2d,8'h2a,8'h24,8'h18,8'h08,8'h00,8'h00,8'h00,8'h00,8'h1b,8'h1e,8'h20,8'h1c,8'h12,8'h12,8'h00,8'h00,8'h00,8'h00,8'h00,8'h11,8'h20,8'h27,8'h24,8'h0f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h37,8'h4d,8'h51,8'h59,8'h4d,8'h00,8'h00,8'h00,8'h1d,8'h2c,8'h32,8'h32,8'h34,8'h34,8'h35,8'h36,8'h35,8'h32,8'h31,8'h32,8'h30,8'h31,8'h34,8'h33,8'h30,8'h2d,8'h2e,8'h30,8'h2f,8'h2f,8'h2d,8'h27,8'h23,8'h1f,8'h1c,8'h00,8'h00,8'h00,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h26,8'h24,8'h00,8'h00,8'h00,8'h11,8'h1f,8'h2b,8'h2d,8'h2f,8'h34,8'h35,8'h37,8'h37,8'h37,8'h37,8'h39,8'h3a,8'h36,8'h37,8'h35,8'h36,8'h37,8'h38,8'h35,8'h33,8'h2f,8'h30,8'h33,8'h35,8'h35,8'h33,8'h33,8'h32,8'h2f,8'h2f,8'h30,8'h2d,8'h38,8'h35,8'h36,8'h38,8'h39,8'h39,8'h3b,8'h3c,8'h39,8'h38,8'h39,8'h36,8'h33,8'h31,8'h34,8'h31,8'h2a,8'h25,8'h17,8'h07,8'h00,8'h00,8'h00,8'h00,8'h0d,8'h21,8'h2d,8'h2f,8'h36,8'h35,8'h3a,8'h38,8'h34,8'h35,8'h36,8'h35,8'h30,8'h2e,8'h2f,8'h31,8'h2d,8'h2b,8'h2d,8'h2d,8'h2f,8'h2e,8'h2b,8'h2c,8'h27,8'h16,8'h00,8'h00,8'h00,8'h00,8'h1e,8'h24,8'h00,8'h00,8'h09,8'h24,8'h2d,8'h30,8'h33,8'h32,8'h32,8'h31,8'h2c,8'h20,8'h00,8'h00,8'h00,8'h22,8'h20,8'h00,8'h00,8'h1f,8'h2f,8'h34,8'h34,8'h31,8'h32,8'h35,8'h33,8'h31,8'h30,8'h2f,8'h31,8'h33,8'h30,8'h2e,8'h2e,8'h2f,8'h2e,8'h30,8'h31,8'h32,8'h30,8'h30,8'h2c,8'h23,8'h12,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1e,8'h28,8'h2a,8'h21,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h29,8'h4d,8'h42,8'h00,8'h00,8'h00,8'h21,8'h2c,8'h2f,8'h33,8'h33,8'h33,8'h34,8'h33,8'h32,8'h33,8'h34,8'h31,8'h30,8'h2f,8'h2f,8'h2c,8'h20,8'h21,8'h30,8'h2f,8'h2e,8'h2b,8'h2a,8'h22,8'h10,8'h0a,8'h00,8'h00,8'h00,8'h24,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h26,8'h24,8'h00,8'h00,8'h00,8'h12,8'h20,8'h28,8'h2c,8'h2f,8'h32,8'h35,8'h36,8'h38,8'h38,8'h38,8'h38,8'h38,8'h39,8'h36,8'h36,8'h37,8'h37,8'h36,8'h35,8'h34,8'h30,8'h35,8'h34,8'h33,8'h33,8'h32,8'h33,8'h31,8'h30,8'h2e,8'h21,8'h1c,8'h36,8'h35,8'h34,8'h35,8'h36,8'h39,8'h3c,8'h3c,8'h34,8'h35,8'h36,8'h32,8'h31,8'h2f,8'h2c,8'h25,8'h22,8'h14,8'h08,8'h00,8'h00,8'h00,8'h00,8'h00,8'h13,8'h21,8'h2f,8'h33,8'h37,8'h38,8'h37,8'h32,8'h33,8'h36,8'h35,8'h32,8'h2e,8'h2d,8'h2d,8'h2a,8'h21,8'h21,8'h2c,8'h2d,8'h2e,8'h2d,8'h29,8'h25,8'h18,8'h02,8'h00,8'h00,8'h00,8'h22,8'h27,8'h25,8'h00,8'h00,8'h0a,8'h24,8'h2c,8'h2f,8'h33,8'h32,8'h31,8'h2e,8'h28,8'h11,8'h00,8'h00,8'h00,8'h22,8'h1b,8'h00,8'h05,8'h22,8'h2b,8'h31,8'h32,8'h30,8'h30,8'h32,8'h32,8'h2f,8'h2f,8'h30,8'h30,8'h32,8'h2e,8'h29,8'h25,8'h23,8'h2d,8'h34,8'h33,8'h33,8'h31,8'h2c,8'h23,8'h10,8'h00,8'h00,8'h00,8'h00,8'h12,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h12,8'h1e,8'h29,8'h2a,8'h20,8'h10,8'h0f,8'h05,8'h0c,8'h18,8'h1e,8'h13,8'h11,8'h14,8'h12,8'h1a,8'h17,8'h11,8'h1a,8'h0d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h1f,8'h00,8'h00,8'h08,8'h21,8'h2c,8'h33,8'h33,8'h34,8'h33,8'h34,8'h30,8'h31,8'h36,8'h34,8'h32,8'h2f,8'h29,8'h24,8'h20,8'h11,8'h1f,8'h2d,8'h2d,8'h2d,8'h28,8'h23,8'h19,8'h15,8'h00,8'h00,8'h00,8'h22,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h26,8'h25,8'h00,8'h00,8'h00,8'h1d,8'h20,8'h28,8'h2b,8'h2c,8'h30,8'h33,8'h34,8'h36,8'h36,8'h39,8'h37,8'h34,8'h36,8'h34,8'h36,8'h37,8'h3b,8'h37,8'h33,8'h32,8'h32,8'h34,8'h33,8'h2f,8'h30,8'h31,8'h2c,8'h29,8'h22,8'h20,8'h0f,8'h1e,8'h35,8'h35,8'h35,8'h34,8'h34,8'h34,8'h36,8'h37,8'h32,8'h30,8'h2f,8'h2b,8'h28,8'h24,8'h1f,8'h1e,8'h0d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h15,8'h23,8'h2e,8'h2f,8'h30,8'h35,8'h32,8'h30,8'h2f,8'h32,8'h31,8'h2f,8'h2c,8'h27,8'h21,8'h1c,8'h1a,8'h1b,8'h26,8'h2d,8'h2c,8'h29,8'h21,8'h1c,8'h01,8'h00,8'h00,8'h00,8'h22,8'h27,8'h27,8'h24,8'h00,8'h00,8'h0f,8'h26,8'h2c,8'h2e,8'h2f,8'h2f,8'h2d,8'h25,8'h1e,8'h0e,8'h00,8'h00,8'h00,8'h24,8'h08,8'h00,8'h1a,8'h26,8'h2e,8'h31,8'h31,8'h31,8'h30,8'h30,8'h2f,8'h2f,8'h31,8'h2d,8'h2d,8'h2a,8'h20,8'h1d,8'h15,8'h18,8'h29,8'h30,8'h2f,8'h2f,8'h2b,8'h24,8'h17,8'h00,8'h00,8'h00,8'h0f,8'h25,8'h25,8'h05,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0c,8'h10,8'h00,8'h00,8'h00,8'h10,8'h1a,8'h25,8'h25,8'h23,8'h1a,8'h12,8'h12,8'h11,8'h16,8'h1f,8'h22,8'h25,8'h2a,8'h2a,8'h29,8'h27,8'h29,8'h28,8'h25,8'h21,8'h21,8'h19,8'h10,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h11,8'h22,8'h2e,8'h31,8'h35,8'h35,8'h33,8'h33,8'h2d,8'h2e,8'h31,8'h2f,8'h2b,8'h23,8'h1d,8'h0f,8'h02,8'h0e,8'h1f,8'h29,8'h2f,8'h2a,8'h23,8'h1d,8'h0f,8'h00,8'h00,8'h00,8'h22,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h26,8'h26,8'h00,8'h00,8'h00,8'h1a,8'h15,8'h27,8'h2b,8'h2b,8'h2f,8'h32,8'h32,8'h32,8'h35,8'h38,8'h35,8'h34,8'h34,8'h35,8'h37,8'h39,8'h39,8'h37,8'h33,8'h32,8'h31,8'h30,8'h30,8'h2f,8'h2d,8'h2c,8'h26,8'h19,8'h09,8'h04,8'h1b,8'h28,8'h32,8'h34,8'h37,8'h35,8'h33,8'h31,8'h32,8'h34,8'h32,8'h2c,8'h28,8'h25,8'h1d,8'h15,8'h0c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h23,8'h26,8'h00,8'h00,8'h12,8'h25,8'h2c,8'h2d,8'h2f,8'h33,8'h32,8'h31,8'h2e,8'h2e,8'h2c,8'h2b,8'h27,8'h20,8'h0a,8'h00,8'h00,8'h11,8'h21,8'h29,8'h28,8'h23,8'h1c,8'h04,8'h00,8'h00,8'h00,8'h23,8'h27,8'h27,8'h27,8'h23,8'h00,8'h00,8'h12,8'h27,8'h2b,8'h2c,8'h2d,8'h2c,8'h28,8'h1f,8'h0f,8'h00,8'h00,8'h00,8'h1f,8'h26,8'h00,8'h00,8'h18,8'h27,8'h30,8'h31,8'h2f,8'h30,8'h30,8'h2f,8'h2e,8'h2c,8'h2e,8'h29,8'h22,8'h19,8'h0f,8'h00,8'h00,8'h14,8'h23,8'h2a,8'h2b,8'h28,8'h20,8'h13,8'h00,8'h00,8'h00,8'h12,8'h26,8'h27,8'h00,8'h25,8'h24,8'h21,8'h23,8'h24,8'h25,8'h26,8'h25,8'h01,8'h00,8'h00,8'h1a,8'h1f,8'h1d,8'h16,8'h13,8'h07,8'h04,8'h09,8'h0c,8'h0d,8'h16,8'h1b,8'h23,8'h2a,8'h30,8'h31,8'h30,8'h30,8'h30,8'h31,8'h2f,8'h2f,8'h28,8'h1f,8'h11,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0f,8'h21,8'h2b,8'h30,8'h32,8'h30,8'h32,8'h30,8'h2d,8'h2b,8'h29,8'h26,8'h1d,8'h16,8'h00,8'h00,8'h00,8'h00,8'h1f,8'h26,8'h2c,8'h24,8'h18,8'h17,8'h00,8'h00,8'h00,8'h23,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h26,8'h07,8'h00,8'h00,8'h0c,8'h15,8'h24,8'h28,8'h2c,8'h30,8'h32,8'h32,8'h33,8'h36,8'h37,8'h36,8'h33,8'h35,8'h36,8'h34,8'h34,8'h32,8'h33,8'h32,8'h30,8'h2e,8'h2c,8'h2d,8'h2b,8'h25,8'h21,8'h1e,8'h00,8'h00,8'h01,8'h1b,8'h29,8'h30,8'h33,8'h34,8'h33,8'h32,8'h31,8'h30,8'h2e,8'h29,8'h23,8'h1c,8'h0e,8'h06,8'h00,8'h00,8'h00,8'h00,8'h00,8'h15,8'h24,8'h27,8'h24,8'h00,8'h00,8'h12,8'h21,8'h2a,8'h2d,8'h2f,8'h32,8'h2f,8'h2e,8'h2c,8'h28,8'h25,8'h20,8'h18,8'h09,8'h00,8'h00,8'h00,8'h14,8'h1f,8'h24,8'h23,8'h12,8'h00,8'h00,8'h00,8'h0a,8'h24,8'h27,8'h27,8'h27,8'h27,8'h24,8'h00,8'h00,8'h19,8'h26,8'h2a,8'h2b,8'h29,8'h24,8'h1a,8'h0c,8'h01,8'h00,8'h00,8'h02,8'h25,8'h26,8'h00,8'h00,8'h17,8'h26,8'h2f,8'h2e,8'h2c,8'h2e,8'h2f,8'h2d,8'h2a,8'h22,8'h22,8'h20,8'h10,8'h00,8'h00,8'h00,8'h00,8'h19,8'h21,8'h26,8'h26,8'h1b,8'h09,8'h00,8'h00,8'h00,8'h1a,8'h26,8'h27,8'h00,8'h00,8'h26,8'h26,8'h26,8'h26,8'h26,8'h26,8'h26,8'h1f,8'h00,8'h00,8'h0f,8'h12,8'h09,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h02,8'h12,8'h17,8'h25,8'h2b,8'h31,8'h33,8'h30,8'h31,8'h32,8'h31,8'h30,8'h2b,8'h23,8'h14,8'h0b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0b,8'h1c,8'h29,8'h2d,8'h2f,8'h2d,8'h29,8'h28,8'h25,8'h20,8'h1f,8'h1e,8'h09,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1e,8'h23,8'h22,8'h13,8'h15,8'h00,8'h00,8'h00,8'h23,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h26,8'h21,8'h00,8'h00,8'h00,8'h1d,8'h1f,8'h24,8'h2c,8'h30,8'h31,8'h31,8'h33,8'h35,8'h35,8'h34,8'h35,8'h35,8'h33,8'h32,8'h32,8'h31,8'h2f,8'h31,8'h2f,8'h29,8'h28,8'h28,8'h22,8'h11,8'h01,8'h00,8'h00,8'h00,8'h0e,8'h1e,8'h2a,8'h32,8'h35,8'h33,8'h31,8'h2e,8'h2e,8'h27,8'h21,8'h18,8'h07,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0b,8'h22,8'h25,8'h26,8'h00,8'h26,8'h23,8'h00,8'h00,8'h11,8'h1a,8'h23,8'h28,8'h2c,8'h2a,8'h27,8'h24,8'h20,8'h17,8'h15,8'h07,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1b,8'h19,8'h15,8'h15,8'h00,8'h00,8'h00,8'h20,8'h26,8'h27,8'h27,8'h27,8'h27,8'h27,8'h24,8'h00,8'h00,8'h19,8'h24,8'h27,8'h26,8'h1f,8'h1a,8'h17,8'h00,8'h00,8'h00,8'h14,8'h25,8'h26,8'h26,8'h11,8'h00,8'h09,8'h21,8'h24,8'h23,8'h22,8'h23,8'h24,8'h21,8'h1e,8'h14,8'h02,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0f,8'h20,8'h23,8'h1b,8'h03,8'h00,8'h00,8'h07,8'h25,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h06,8'h12,8'h24,8'h2e,8'h33,8'h32,8'h31,8'h32,8'h33,8'h36,8'h32,8'h2f,8'h27,8'h17,8'h0c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h19,8'h21,8'h21,8'h21,8'h21,8'h1a,8'h18,8'h0d,8'h0b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h12,8'h18,8'h15,8'h12,8'h00,8'h00,8'h00,8'h24,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h26,8'h26,8'h04,8'h00,8'h00,8'h13,8'h16,8'h20,8'h26,8'h2d,8'h2f,8'h31,8'h32,8'h34,8'h34,8'h35,8'h34,8'h33,8'h32,8'h30,8'h30,8'h30,8'h30,8'h2f,8'h2c,8'h29,8'h23,8'h1a,8'h0a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h19,8'h21,8'h2d,8'h30,8'h30,8'h2c,8'h2a,8'h25,8'h21,8'h12,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h21,8'h26,8'h26,8'h26,8'h00,8'h00,8'h26,8'h24,8'h00,8'h00,8'h00,8'h16,8'h16,8'h1b,8'h1f,8'h1b,8'h1b,8'h1a,8'h0d,8'h01,8'h00,8'h00,8'h00,8'h00,8'h14,8'h00,8'h00,8'h09,8'h14,8'h07,8'h00,8'h00,8'h00,8'h17,8'h26,8'h00,8'h27,8'h27,8'h27,8'h27,8'h27,8'h24,8'h00,8'h00,8'h16,8'h18,8'h20,8'h18,8'h10,8'h15,8'h00,8'h00,8'h00,8'h1a,8'h26,8'h26,8'h00,8'h26,8'h22,8'h00,8'h00,8'h20,8'h1b,8'h10,8'h0d,8'h15,8'h15,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h21,8'h19,8'h00,8'h00,8'h18,8'h1d,8'h0b,8'h00,8'h00,8'h00,8'h26,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0b,8'h06,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'h17,8'h27,8'h30,8'h30,8'h32,8'h35,8'h34,8'h34,8'h33,8'h34,8'h30,8'h24,8'h1f,8'h04,8'h00,8'h00,8'h00,8'h00,8'h05,8'h1d,8'h15,8'h10,8'h0b,8'h0c,8'h11,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1f,8'h00,8'h00,8'h00,8'h1f,8'h15,8'h0f,8'h00,8'h00,8'h00,8'h23,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h26,8'h1d,8'h00,8'h00,8'h04,8'h16,8'h18,8'h21,8'h28,8'h2e,8'h2e,8'h2d,8'h2f,8'h32,8'h31,8'h31,8'h31,8'h2e,8'h2c,8'h2d,8'h2e,8'h2b,8'h26,8'h23,8'h23,8'h0e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h15,8'h23,8'h2b,8'h2d,8'h2b,8'h24,8'h1d,8'h1e,8'h0d,8'h0a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h1f,8'h00,8'h00,8'h00,8'h1f,8'h15,8'h0e,8'h08,8'h07,8'h00,8'h00,8'h00,8'h00,8'h00,8'h09,8'h24,8'h26,8'h1b,8'h00,8'h00,8'h19,8'h00,8'h00,8'h00,8'h1f,8'h26,8'h26,8'h00,8'h27,8'h27,8'h27,8'h27,8'h27,8'h24,8'h00,8'h00,8'h15,8'h0c,8'h15,8'h15,8'h00,8'h00,8'h00,8'h00,8'h21,8'h27,8'h27,8'h00,8'h00,8'h26,8'h25,8'h02,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h12,8'h22,8'h27,8'h27,8'h23,8'h00,8'h00,8'h16,8'h07,8'h00,8'h00,8'h00,8'h24,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h25,8'h00,8'h00,8'h00,8'h00,8'h11,8'h21,8'h25,8'h26,8'h26,8'h23,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0e,8'h22,8'h2c,8'h2f,8'h34,8'h37,8'h36,8'h32,8'h33,8'h35,8'h2f,8'h27,8'h23,8'h13,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h23,8'h26,8'h26,8'h16,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h21,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h26,8'h25,8'h00,8'h00,8'h00,8'h14,8'h1b,8'h1b,8'h20,8'h2a,8'h2a,8'h29,8'h2b,8'h2c,8'h2e,8'h2f,8'h2f,8'h2d,8'h2b,8'h28,8'h25,8'h1b,8'h11,8'h0f,8'h0c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h10,8'h17,8'h27,8'h2d,8'h28,8'h1f,8'h14,8'h12,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h21,8'h26,8'h00,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h18,8'h23,8'h26,8'h26,8'h00,8'h1f,8'h00,8'h00,8'h00,8'h00,8'h00,8'h23,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h27,8'h26,8'h06,8'h00,8'h00,8'h10,8'h12,8'h00,8'h00,8'h00,8'h05,8'h23,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h06,8'h1f,8'h25,8'h27,8'h00,8'h27,8'h27,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h08,8'h25,8'h27,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h22,8'h00,8'h06,8'h22,8'h26,8'h26,8'h00,8'h26,8'h26,8'h26,8'h0d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h16,8'h27,8'h2f,8'h33,8'h36,8'h34,8'h33,8'h31,8'h34,8'h31,8'h2a,8'h23,8'h0e,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1b,8'h23,8'h26,8'h00,8'h26,8'h00,8'h26,8'h0d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h17,8'h00,8'h00,8'h00,8'h07,8'h16,8'h15,8'h1f,8'h1c,8'h1e,8'h21,8'h24,8'h29,8'h26,8'h25,8'h25,8'h22,8'h20,8'h1e,8'h17,8'h06,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1a,8'h1d,8'h25,8'h23,8'h1f,8'h0c,8'h08,8'h00,8'h00,8'h00,8'h00,8'h00,8'h13,8'h24,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0c,8'h21,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h16,8'h00,8'h00,8'h00,8'h24,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h27,8'h22,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h20,8'h00,8'h00,8'h00,8'h15,8'h20,8'h22,8'h25,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h10,8'h00,8'h00,8'h00,8'h07,8'h25,8'h27,8'h27,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h24,8'h22,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h0f,8'h00,8'h00,8'h00,8'h09,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h11,8'h22,8'h2e,8'h33,8'h35,8'h34,8'h34,8'h33,8'h34,8'h32,8'h2e,8'h26,8'h11,8'h00,8'h00,8'h00,8'h07,8'h22,8'h0b,8'h00,8'h00,8'h00,8'h0b,8'h20,8'h25,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h13,8'h01,8'h00,8'h0c,8'h23,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h26,8'h1a,8'h00,8'h00,8'h00,8'h00,8'h10,8'h20,8'h1b,8'h12,8'h11,8'h18,8'h1d,8'h17,8'h15,8'h0f,8'h10,8'h16,8'h1f,8'h08,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h19,8'h00,8'h00,8'h00,8'h14,8'h15,8'h1e,8'h09,8'h07,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1f,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h25,8'h24,8'h25,8'h25,8'h24,8'h24,8'h25,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h25,8'h24,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h27,8'h27,8'h27,8'h26,8'h1a,8'h00,8'h00,8'h00,8'h00,8'h23,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h25,8'h25,8'h26,8'h00,8'h26,8'h26,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h1a,8'h1b,8'h23,8'h25,8'h26,8'h00,8'h27,8'h27,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h1a,8'h00,8'h00,8'h00,8'h0e,8'h0a,8'h00,8'h00,8'h00,8'h00,8'h24,8'h0e,8'h00,8'h00,8'h0b,8'h1e,8'h2b,8'h31,8'h34,8'h35,8'h35,8'h34,8'h32,8'h33,8'h30,8'h27,8'h10,8'h00,8'h00,8'h00,8'h10,8'h26,8'h25,8'h25,8'h26,8'h25,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h25,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h21,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h09,8'h0a,8'h06,8'h02,8'h0b,8'h07,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h15,8'h24,8'h25,8'h25,8'h00,8'h00,8'h10,8'h11,8'h0e,8'h0b,8'h00,8'h00,8'h00,8'h00,8'h00,8'h20,8'h25,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h26,8'h26,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h25,8'h24,8'h24,8'h25,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h25,8'h1c,8'h00,8'h00,8'h00,8'h0f,8'h12,8'h03,8'h00,8'h00,8'h00,8'h21,8'h27,8'h21,8'h00,8'h00,8'h07,8'h15,8'h28,8'h31,8'h35,8'h35,8'h36,8'h35,8'h34,8'h33,8'h30,8'h28,8'h15,8'h00,8'h00,8'h00,8'h21,8'h00,8'h26,8'h26,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h10,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0e,8'h23,8'h26,8'h26,8'h26,8'h22,8'h00,8'h00,8'h13,8'h12,8'h00,8'h00,8'h00,8'h00,8'h00,8'h17,8'h25,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h17,8'h00,8'h00,8'h00,8'h16,8'h0e,8'h0a,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h20,8'h00,8'h00,8'h00,8'h0e,8'h27,8'h30,8'h34,8'h33,8'h35,8'h34,8'h35,8'h33,8'h2d,8'h24,8'h14,8'h00,8'h00,8'h00,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h1e,8'h09,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h15,8'h25,8'h26,8'h00,8'h00,8'h00,8'h00,8'h15,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h18,8'h22,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h19,8'h00,8'h00,8'h00,8'h09,8'h0f,8'h12,8'h03,8'h00,8'h00,8'h00,8'h21,8'h24,8'h13,8'h00,8'h00,8'h00,8'h09,8'h15,8'h2a,8'h2d,8'h2f,8'h32,8'h32,8'h32,8'h32,8'h30,8'h2b,8'h20,8'h13,8'h00,8'h00,8'h1a,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h23,8'h22,8'h20,8'h19,8'h19,8'h17,8'h1e,8'h23,8'h24,8'h25,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h26,8'h04,8'h00,8'h00,8'h00,8'h00,8'h02,8'h24,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h17,8'h00,8'h00,8'h00,8'h17,8'h1c,8'h19,8'h0e,8'h00,8'h00,8'h00,8'h05,8'h22,8'h00,8'h00,8'h00,8'h00,8'h0e,8'h17,8'h26,8'h2e,8'h31,8'h32,8'h33,8'h30,8'h31,8'h31,8'h2d,8'h25,8'h13,8'h0a,8'h00,8'h00,8'h23,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h26,8'h26,8'h26,8'h00,8'h26,8'h00,8'h26,8'h26,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h00,8'h00,8'h00,8'h00,8'h1f,8'h25,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h27,8'h22,8'h00,8'h00,8'h00,8'h10,8'h1a,8'h21,8'h18,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0f,8'h19,8'h26,8'h2d,8'h30,8'h32,8'h33,8'h33,8'h32,8'h31,8'h30,8'h2a,8'h21,8'h0f,8'h00,8'h00,8'h00,8'h25,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h21,8'h00,8'h18,8'h24,8'h26,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h1e,8'h00,8'h00,8'h00,8'h14,8'h20,8'h23,8'h22,8'h0a,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h08,8'h17,8'h1f,8'h28,8'h2c,8'h31,8'h33,8'h31,8'h31,8'h31,8'h2f,8'h2e,8'h2d,8'h22,8'h10,8'h02,8'h00,8'h00,8'h1a,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h24,8'h0c,8'h00,8'h00,8'h04,8'h13,8'h19,8'h24,8'h21,8'h14,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0c,8'h15,8'h21,8'h29,8'h2f,8'h2f,8'h30,8'h32,8'h31,8'h30,8'h2f,8'h2c,8'h28,8'h26,8'h14,8'h08,8'h00,8'h00,8'h00,8'h24,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h00,8'h00,8'h00,8'h00,8'h16,8'h19,8'h22,8'h23,8'h16,8'h09,8'h00,8'h00,8'h00,8'h00,8'h00,8'h05,8'h16,8'h1a,8'h25,8'h2b,8'h2f,8'h30,8'h31,8'h30,8'h30,8'h32,8'h31,8'h2e,8'h2a,8'h24,8'h1e,8'h18,8'h00,8'h00,8'h00,8'h20,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h1f,8'h00,8'h00,8'h00,8'h10,8'h16,8'h20,8'h25,8'h26,8'h20,8'h08,8'h00,8'h00,8'h00,8'h00,8'h00,8'h10,8'h18,8'h25,8'h28,8'h2c,8'h2e,8'h2e,8'h30,8'h31,8'h30,8'h2f,8'h2f,8'h2d,8'h2b,8'h26,8'h19,8'h13,8'h00,8'h00,8'h00,8'h1d,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h1f,8'h00,8'h00,8'h00,8'h10,8'h19,8'h1e,8'h26,8'h2a,8'h27,8'h1a,8'h00,8'h00,8'h00,8'h00,8'h07,8'h16,8'h1e,8'h26,8'h2b,8'h2a,8'h2d,8'h2f,8'h2e,8'h2f,8'h2e,8'h2f,8'h2f,8'h2b,8'h28,8'h23,8'h1a,8'h0d,8'h00,8'h00,8'h00,8'h09,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h1e,8'h00,8'h00,8'h00,8'h11,8'h13,8'h20,8'h24,8'h27,8'h29,8'h21,8'h0f,8'h00,8'h00,8'h0b,8'h11,8'h1a,8'h22,8'h29,8'h2c,8'h2c,8'h2d,8'h2f,8'h2e,8'h2f,8'h2e,8'h2e,8'h2e,8'h2e,8'h27,8'h21,8'h18,8'h0d,8'h00,8'h00,8'h00,8'h00,8'h24,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h17,8'h00,8'h00,8'h1b,8'h13,8'h1f,8'h25,8'h26,8'h27,8'h29,8'h17,8'h0a,8'h0c,8'h12,8'h1f,8'h23,8'h28,8'h2c,8'h2d,8'h2e,8'h2d,8'h2c,8'h2e,8'h2f,8'h2f,8'h2f,8'h2c,8'h2c,8'h2a,8'h21,8'h13,8'h00,8'h00,8'h00,8'h00,8'h14,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h1f,8'h00,8'h00,8'h10,8'h1c,8'h25,8'h29,8'h2b,8'h2a,8'h2b,8'h24,8'h1a,8'h20,8'h26,8'h2a,8'h2c,8'h2b,8'h2f,8'h30,8'h2f,8'h2e,8'h2d,8'h30,8'h2f,8'h2e,8'h2d,8'h29,8'h28,8'h22,8'h11,8'h04,8'h00,8'h00,8'h00,8'h19,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h20,8'h00,8'h00,8'h0d,8'h17,8'h24,8'h2a,8'h2c,8'h2b,8'h2c,8'h2c,8'h2b,8'h2b,8'h2d,8'h2f,8'h31,8'h30,8'h2f,8'h2f,8'h2e,8'h2e,8'h2f,8'h2e,8'h2c,8'h2c,8'h29,8'h23,8'h1d,8'h1b,8'h00,8'h00,8'h00,8'h00,8'h1e,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h20,8'h00,8'h00,8'h07,8'h13,8'h25,8'h2b,8'h2b,8'h2b,8'h2d,8'h2d,8'h2e,8'h2b,8'h2b,8'h2e,8'h2e,8'h2e,8'h2e,8'h2f,8'h2e,8'h2e,8'h2e,8'h2c,8'h28,8'h27,8'h27,8'h18,8'h09,8'h00,8'h00,8'h00,8'h00,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h22,8'h00,8'h00,8'h06,8'h11,8'h23,8'h2a,8'h2c,8'h2a,8'h2c,8'h2f,8'h30,8'h2d,8'h2e,8'h2f,8'h2e,8'h2d,8'h2e,8'h2e,8'h2d,8'h2c,8'h2e,8'h29,8'h24,8'h1e,8'h19,8'h01,8'h00,8'h00,8'h00,8'h00,8'h23,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h25,8'h00,8'h00,8'h00,8'h12,8'h23,8'h29,8'h2b,8'h2b,8'h2c,8'h2f,8'h30,8'h2e,8'h2f,8'h30,8'h2f,8'h2d,8'h2b,8'h2c,8'h2c,8'h2a,8'h29,8'h24,8'h1f,8'h11,8'h00,8'h00,8'h00,8'h00,8'h03,8'h24,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h25,8'h00,8'h00,8'h00,8'h12,8'h25,8'h29,8'h29,8'h2a,8'h2d,8'h2c,8'h2c,8'h2c,8'h2e,8'h2f,8'h2d,8'h2c,8'h2a,8'h2a,8'h29,8'h26,8'h22,8'h18,8'h06,8'h00,8'h00,8'h00,8'h00,8'h1b,8'h25,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h25,8'h00,8'h00,8'h00,8'h17,8'h25,8'h27,8'h29,8'h2a,8'h2c,8'h2b,8'h2c,8'h2d,8'h2d,8'h2e,8'h2b,8'h2a,8'h27,8'h27,8'h24,8'h1f,8'h16,8'h02,8'h00,8'h00,8'h00,8'h00,8'h1f,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h00,8'h00,8'h00,8'h17,8'h24,8'h26,8'h29,8'h28,8'h2b,8'h2b,8'h2c,8'h2c,8'h2d,8'h2d,8'h2a,8'h26,8'h24,8'h23,8'h1e,8'h16,8'h09,8'h00,8'h00,8'h00,8'h00,8'h22,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h00,8'h00,8'h00,8'h12,8'h22,8'h25,8'h29,8'h27,8'h2b,8'h2b,8'h2b,8'h2b,8'h2a,8'h2b,8'h2a,8'h26,8'h24,8'h1e,8'h0c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h09,8'h00,8'h00,8'h12,8'h1c,8'h26,8'h28,8'h27,8'h2a,8'h2b,8'h2a,8'h29,8'h27,8'h26,8'h23,8'h21,8'h15,8'h06,8'h00,8'h00,8'h00,8'h00,8'h03,8'h23,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h09,8'h00,8'h00,8'h13,8'h19,8'h24,8'h26,8'h27,8'h2a,8'h29,8'h27,8'h25,8'h24,8'h20,8'h14,8'h0d,8'h00,8'h00,8'h00,8'h00,8'h01,8'h24,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h09,8'h00,8'h00,8'h0e,8'h14,8'h22,8'h25,8'h26,8'h27,8'h26,8'h23,8'h20,8'h17,8'h17,8'h05,8'h00,8'h00,8'h00,8'h00,8'h12,8'h25,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h10,8'h00,8'h00,8'h0c,8'h14,8'h24,8'h24,8'h25,8'h23,8'h21,8'h1a,8'h15,8'h10,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1f,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0e,8'h00,8'h00,8'h14,8'h1a,8'h23,8'h22,8'h21,8'h21,8'h16,8'h0d,8'h00,8'h00,8'h00,8'h00,8'h00,8'h15,8'h25,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0d,8'h00,8'h00,8'h19,8'h1f,8'h22,8'h24,8'h1d,8'h0f,8'h03,8'h00,8'h00,8'h00,8'h00,8'h00,8'h1f,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0d,8'h00,8'h00,8'h13,8'h10,8'h1d,8'h1e,8'h17,8'h00,8'h00,8'h00,8'h00,8'h00,8'h03,8'h24,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h09,8'h00,8'h00,8'h12,8'h0e,8'h0c,8'h00,8'h00,8'h00,8'h00,8'h00,8'h08,8'h25,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h00,8'h00,8'h17,8'h07,8'h00,8'h00,8'h00,8'h00,8'h00,8'h12,8'h25,8'h00,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h09,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h0f,8'h23,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h08,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h22,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h25,8'h00,8'h00,8'h00,8'h00,8'h00,8'h06,8'h23,8'h00,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h24,8'h00,8'h00,8'h00,8'h12,8'h21,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h00,8'h00,8'h23,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h24,8'h26,8'h27,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},
'{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h26,8'h26,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}};

assign SpriteR = SpriteTableR[SpriteY][SpriteX];
assign SpriteG = SpriteTableG[SpriteY][SpriteX];
assign SpriteB = SpriteTableB[SpriteY][SpriteX];

endmodule
